`timescale 1ns / 1ps
`include "cnu.v"
`include "vnu.v"
`include "vnu_1.v"
`include "vnu_h.v"
module decode(clk, rst, data_0 ,data_1 ,data_2 ,data_3 ,data_4 ,data_5 ,data_6 ,data_7 ,data_8 ,data_9 ,data_10 ,data_11 ,data_12 ,data_13 ,data_14 ,data_15 ,data_16 ,data_17 ,data_18 ,data_19 ,data_20 ,data_21 ,data_22 ,data_23 ,data_24 ,data_25 ,data_26 ,data_27 ,data_28 ,data_29 ,data_30 ,data_31 ,data_32 ,data_33 ,data_34 ,data_35 ,data_36 ,data_37 ,data_38 ,data_39 ,data_40 ,data_41 ,data_42 ,data_43 ,data_44 ,data_45 ,data_46 ,data_47 ,data_48 ,data_49 ,data_50 ,data_51 ,data_52 ,data_53 ,data_54 ,data_55 ,data_56 ,data_57 ,data_58 ,data_59 ,data_60 ,data_61 ,data_62 ,data_63 ,data_64 ,data_65 ,data_66 ,data_67 ,data_68 ,data_69 ,data_70 ,data_71 ,data_72 ,data_73 ,data_74 ,data_75 ,data_76 ,data_77 ,data_78 ,data_79 ,data_80 ,data_81 ,data_82 ,data_83 ,data_84 ,data_85 ,data_86 ,data_87 ,data_88 ,data_89 ,data_90 ,data_91 ,data_92 ,data_93 ,data_94 ,data_95 ,data_96 ,data_97 ,data_98 ,data_99 ,data_100 ,data_101 ,data_102 ,data_103 ,data_104 ,data_105 ,data_106 ,data_107 ,data_108 ,data_109 ,data_110 ,data_111 ,data_112 ,data_113 ,data_114 ,data_115 ,data_116 ,data_117 ,data_118 ,data_119 ,data_120 ,data_121 ,data_122 ,data_123 ,data_124 ,data_125 ,data_126 ,data_127 ,data_128 ,data_129 ,data_130 ,data_131 ,data_132 ,data_133 ,data_134 ,data_135 ,data_136 ,data_137 ,data_138 ,data_139 ,data_140 ,data_141 ,data_142 ,data_143 ,data_144 ,data_145 ,data_146 ,data_147 ,data_148 ,data_149 ,data_150 ,data_151 ,data_152 ,data_153 ,data_154 ,data_155 ,data_156 ,data_157 ,data_158 ,data_159 ,data_160 ,data_161 ,data_162 ,data_163 ,data_164 ,data_165 ,data_166 ,data_167 ,data_168 ,data_169 ,data_170 ,data_171 ,data_172 ,data_173 ,data_174 ,data_175 ,data_176 ,data_177 ,data_178 ,data_179 ,data_180 ,data_181 ,data_182 ,data_183 ,data_184 ,data_185 ,data_186 ,data_187 ,data_188 ,data_189 ,data_190 ,data_191 ,data_192 ,data_193 ,data_194 ,data_195 ,data_196 ,data_197, data_out);

//receive input data of 5*211 size. send repective data to all bit nodes as intrinsic info. receive corresponding bit to check msgs from bit nodes. send correct bit to check msgs to check nodes and receive chk to bit msgs. repeat for 15 iterations and then perform hard decoding. 

input [7:0] data_0 ,data_1 ,data_2 ,data_3 ,data_4 ,data_5 ,data_6 ,data_7 ,data_8 ,data_9 ,data_10 ,data_11 ,data_12 ,data_13 ,data_14 ,data_15 ,data_16 ,data_17 ,data_18 ,data_19 ,data_20 ,data_21 ,data_22 ,data_23 ,data_24 ,data_25 ,data_26 ,data_27 ,data_28 ,data_29 ,data_30 ,data_31 ,data_32 ,data_33 ,data_34 ,data_35 ,data_36 ,data_37 ,data_38 ,data_39 ,data_40 ,data_41 ,data_42 ,data_43 ,data_44 ,data_45 ,data_46 ,data_47 ,data_48 ,data_49 ,data_50 ,data_51 ,data_52 ,data_53 ,data_54 ,data_55 ,data_56 ,data_57 ,data_58 ,data_59 ,data_60 ,data_61 ,data_62 ,data_63 ,data_64 ,data_65 ,data_66 ,data_67 ,data_68 ,data_69 ,data_70 ,data_71 ,data_72 ,data_73 ,data_74 ,data_75 ,data_76 ,data_77 ,data_78 ,data_79 ,data_80 ,data_81 ,data_82 ,data_83 ,data_84 ,data_85 ,data_86 ,data_87 ,data_88 ,data_89 ,data_90 ,data_91 ,data_92 ,data_93 ,data_94 ,data_95 ,data_96 ,data_97 ,data_98 ,data_99 ,data_100 ,data_101 ,data_102 ,data_103 ,data_104 ,data_105 ,data_106 ,data_107 ,data_108 ,data_109 ,data_110 ,data_111 ,data_112 ,data_113 ,data_114 ,data_115 ,data_116 ,data_117 ,data_118 ,data_119 ,data_120 ,data_121 ,data_122 ,data_123 ,data_124 ,data_125 ,data_126 ,data_127 ,data_128 ,data_129 ,data_130 ,data_131 ,data_132 ,data_133 ,data_134 ,data_135 ,data_136 ,data_137 ,data_138 ,data_139 ,data_140 ,data_141 ,data_142 ,data_143 ,data_144 ,data_145 ,data_146 ,data_147 ,data_148 ,data_149 ,data_150 ,data_151 ,data_152 ,data_153 ,data_154 ,data_155 ,data_156 ,data_157 ,data_158 ,data_159 ,data_160 ,data_161 ,data_162 ,data_163 ,data_164 ,data_165 ,data_166 ,data_167 ,data_168 ,data_169 ,data_170 ,data_171 ,data_172 ,data_173 ,data_174 ,data_175 ,data_176 ,data_177 ,data_178 ,data_179 ,data_180 ,data_181 ,data_182 ,data_183 ,data_184 ,data_185 ,data_186 ,data_187 ,data_188 ,data_189 ,data_190 ,data_191 ,data_192 ,data_193 ,data_194 ,data_195 ,data_196 ,data_197;
input clk, rst;
output [0:197]data_out;
//input data_in_en;
wire [7:0] msg_to_check_it_0_cnu_0_in_0, msg_to_check_it_0_cnu_0_in_1, msg_to_check_it_0_cnu_0_in_2, msg_to_check_it_0_cnu_0_in_3, msg_to_check_it_0_cnu_0_in_4, msg_to_check_it_0_cnu_0_in_5, msg_to_check_it_0_cnu_1_in_0, msg_to_check_it_0_cnu_1_in_1, msg_to_check_it_0_cnu_1_in_2, msg_to_check_it_0_cnu_1_in_3, msg_to_check_it_0_cnu_1_in_4, msg_to_check_it_0_cnu_1_in_5, msg_to_check_it_0_cnu_2_in_0, msg_to_check_it_0_cnu_2_in_1, msg_to_check_it_0_cnu_2_in_2, msg_to_check_it_0_cnu_2_in_3, msg_to_check_it_0_cnu_2_in_4, msg_to_check_it_0_cnu_2_in_5, msg_to_check_it_0_cnu_3_in_0, msg_to_check_it_0_cnu_3_in_1, msg_to_check_it_0_cnu_3_in_2, msg_to_check_it_0_cnu_3_in_3, msg_to_check_it_0_cnu_3_in_4, msg_to_check_it_0_cnu_3_in_5, msg_to_check_it_0_cnu_4_in_0, msg_to_check_it_0_cnu_4_in_1, msg_to_check_it_0_cnu_4_in_2, msg_to_check_it_0_cnu_4_in_3, msg_to_check_it_0_cnu_4_in_4, msg_to_check_it_0_cnu_4_in_5, msg_to_check_it_0_cnu_5_in_0, msg_to_check_it_0_cnu_5_in_1, msg_to_check_it_0_cnu_5_in_2, msg_to_check_it_0_cnu_5_in_3, msg_to_check_it_0_cnu_5_in_4, msg_to_check_it_0_cnu_5_in_5, msg_to_check_it_0_cnu_6_in_0, msg_to_check_it_0_cnu_6_in_1, msg_to_check_it_0_cnu_6_in_2, msg_to_check_it_0_cnu_6_in_3, msg_to_check_it_0_cnu_6_in_4, msg_to_check_it_0_cnu_6_in_5, msg_to_check_it_0_cnu_7_in_0, msg_to_check_it_0_cnu_7_in_1, msg_to_check_it_0_cnu_7_in_2, msg_to_check_it_0_cnu_7_in_3, msg_to_check_it_0_cnu_7_in_4, msg_to_check_it_0_cnu_7_in_5, msg_to_check_it_0_cnu_8_in_0, msg_to_check_it_0_cnu_8_in_1, msg_to_check_it_0_cnu_8_in_2, msg_to_check_it_0_cnu_8_in_3, msg_to_check_it_0_cnu_8_in_4, msg_to_check_it_0_cnu_8_in_5, msg_to_check_it_0_cnu_9_in_0, msg_to_check_it_0_cnu_9_in_1, msg_to_check_it_0_cnu_9_in_2, msg_to_check_it_0_cnu_9_in_3, msg_to_check_it_0_cnu_9_in_4, msg_to_check_it_0_cnu_9_in_5, msg_to_check_it_0_cnu_10_in_0, msg_to_check_it_0_cnu_10_in_1, msg_to_check_it_0_cnu_10_in_2, msg_to_check_it_0_cnu_10_in_3, msg_to_check_it_0_cnu_10_in_4, msg_to_check_it_0_cnu_10_in_5, msg_to_check_it_0_cnu_11_in_0, msg_to_check_it_0_cnu_11_in_1, msg_to_check_it_0_cnu_11_in_2, msg_to_check_it_0_cnu_11_in_3, msg_to_check_it_0_cnu_11_in_4, msg_to_check_it_0_cnu_11_in_5, msg_to_check_it_0_cnu_12_in_0, msg_to_check_it_0_cnu_12_in_1, msg_to_check_it_0_cnu_12_in_2, msg_to_check_it_0_cnu_12_in_3, msg_to_check_it_0_cnu_12_in_4, msg_to_check_it_0_cnu_12_in_5, msg_to_check_it_0_cnu_13_in_0, msg_to_check_it_0_cnu_13_in_1, msg_to_check_it_0_cnu_13_in_2, msg_to_check_it_0_cnu_13_in_3, msg_to_check_it_0_cnu_13_in_4, msg_to_check_it_0_cnu_13_in_5, msg_to_check_it_0_cnu_14_in_0, msg_to_check_it_0_cnu_14_in_1, msg_to_check_it_0_cnu_14_in_2, msg_to_check_it_0_cnu_14_in_3, msg_to_check_it_0_cnu_14_in_4, msg_to_check_it_0_cnu_14_in_5, msg_to_check_it_0_cnu_15_in_0, msg_to_check_it_0_cnu_15_in_1, msg_to_check_it_0_cnu_15_in_2, msg_to_check_it_0_cnu_15_in_3, msg_to_check_it_0_cnu_15_in_4, msg_to_check_it_0_cnu_15_in_5, msg_to_check_it_0_cnu_16_in_0, msg_to_check_it_0_cnu_16_in_1, msg_to_check_it_0_cnu_16_in_2, msg_to_check_it_0_cnu_16_in_3, msg_to_check_it_0_cnu_16_in_4, msg_to_check_it_0_cnu_16_in_5, msg_to_check_it_0_cnu_17_in_0, msg_to_check_it_0_cnu_17_in_1, msg_to_check_it_0_cnu_17_in_2, msg_to_check_it_0_cnu_17_in_3, msg_to_check_it_0_cnu_17_in_4, msg_to_check_it_0_cnu_17_in_5, msg_to_check_it_0_cnu_18_in_0, msg_to_check_it_0_cnu_18_in_1, msg_to_check_it_0_cnu_18_in_2, msg_to_check_it_0_cnu_18_in_3, msg_to_check_it_0_cnu_18_in_4, msg_to_check_it_0_cnu_18_in_5, msg_to_check_it_0_cnu_19_in_0, msg_to_check_it_0_cnu_19_in_1, msg_to_check_it_0_cnu_19_in_2, msg_to_check_it_0_cnu_19_in_3, msg_to_check_it_0_cnu_19_in_4, msg_to_check_it_0_cnu_19_in_5, msg_to_check_it_0_cnu_20_in_0, msg_to_check_it_0_cnu_20_in_1, msg_to_check_it_0_cnu_20_in_2, msg_to_check_it_0_cnu_20_in_3, msg_to_check_it_0_cnu_20_in_4, msg_to_check_it_0_cnu_20_in_5, msg_to_check_it_0_cnu_21_in_0, msg_to_check_it_0_cnu_21_in_1, msg_to_check_it_0_cnu_21_in_2, msg_to_check_it_0_cnu_21_in_3, msg_to_check_it_0_cnu_21_in_4, msg_to_check_it_0_cnu_21_in_5, msg_to_check_it_0_cnu_22_in_0, msg_to_check_it_0_cnu_22_in_1, msg_to_check_it_0_cnu_22_in_2, msg_to_check_it_0_cnu_22_in_3, msg_to_check_it_0_cnu_22_in_4, msg_to_check_it_0_cnu_22_in_5, msg_to_check_it_0_cnu_23_in_0, msg_to_check_it_0_cnu_23_in_1, msg_to_check_it_0_cnu_23_in_2, msg_to_check_it_0_cnu_23_in_3, msg_to_check_it_0_cnu_23_in_4, msg_to_check_it_0_cnu_23_in_5, msg_to_check_it_0_cnu_24_in_0, msg_to_check_it_0_cnu_24_in_1, msg_to_check_it_0_cnu_24_in_2, msg_to_check_it_0_cnu_24_in_3, msg_to_check_it_0_cnu_24_in_4, msg_to_check_it_0_cnu_24_in_5, msg_to_check_it_0_cnu_25_in_0, msg_to_check_it_0_cnu_25_in_1, msg_to_check_it_0_cnu_25_in_2, msg_to_check_it_0_cnu_25_in_3, msg_to_check_it_0_cnu_25_in_4, msg_to_check_it_0_cnu_25_in_5, msg_to_check_it_0_cnu_26_in_0, msg_to_check_it_0_cnu_26_in_1, msg_to_check_it_0_cnu_26_in_2, msg_to_check_it_0_cnu_26_in_3, msg_to_check_it_0_cnu_26_in_4, msg_to_check_it_0_cnu_26_in_5, msg_to_check_it_0_cnu_27_in_0, msg_to_check_it_0_cnu_27_in_1, msg_to_check_it_0_cnu_27_in_2, msg_to_check_it_0_cnu_27_in_3, msg_to_check_it_0_cnu_27_in_4, msg_to_check_it_0_cnu_27_in_5, msg_to_check_it_0_cnu_28_in_0, msg_to_check_it_0_cnu_28_in_1, msg_to_check_it_0_cnu_28_in_2, msg_to_check_it_0_cnu_28_in_3, msg_to_check_it_0_cnu_28_in_4, msg_to_check_it_0_cnu_28_in_5, msg_to_check_it_0_cnu_29_in_0, msg_to_check_it_0_cnu_29_in_1, msg_to_check_it_0_cnu_29_in_2, msg_to_check_it_0_cnu_29_in_3, msg_to_check_it_0_cnu_29_in_4, msg_to_check_it_0_cnu_29_in_5, msg_to_check_it_0_cnu_30_in_0, msg_to_check_it_0_cnu_30_in_1, msg_to_check_it_0_cnu_30_in_2, msg_to_check_it_0_cnu_30_in_3, msg_to_check_it_0_cnu_30_in_4, msg_to_check_it_0_cnu_30_in_5, msg_to_check_it_0_cnu_31_in_0, msg_to_check_it_0_cnu_31_in_1, msg_to_check_it_0_cnu_31_in_2, msg_to_check_it_0_cnu_31_in_3, msg_to_check_it_0_cnu_31_in_4, msg_to_check_it_0_cnu_31_in_5, msg_to_check_it_0_cnu_32_in_0, msg_to_check_it_0_cnu_32_in_1, msg_to_check_it_0_cnu_32_in_2, msg_to_check_it_0_cnu_32_in_3, msg_to_check_it_0_cnu_32_in_4, msg_to_check_it_0_cnu_32_in_5, msg_to_check_it_0_cnu_33_in_0, msg_to_check_it_0_cnu_33_in_1, msg_to_check_it_0_cnu_33_in_2, msg_to_check_it_0_cnu_33_in_3, msg_to_check_it_0_cnu_33_in_4, msg_to_check_it_0_cnu_33_in_5, msg_to_check_it_0_cnu_34_in_0, msg_to_check_it_0_cnu_34_in_1, msg_to_check_it_0_cnu_34_in_2, msg_to_check_it_0_cnu_34_in_3, msg_to_check_it_0_cnu_34_in_4, msg_to_check_it_0_cnu_34_in_5, msg_to_check_it_0_cnu_35_in_0, msg_to_check_it_0_cnu_35_in_1, msg_to_check_it_0_cnu_35_in_2, msg_to_check_it_0_cnu_35_in_3, msg_to_check_it_0_cnu_35_in_4, msg_to_check_it_0_cnu_35_in_5, msg_to_check_it_0_cnu_36_in_0, msg_to_check_it_0_cnu_36_in_1, msg_to_check_it_0_cnu_36_in_2, msg_to_check_it_0_cnu_36_in_3, msg_to_check_it_0_cnu_36_in_4, msg_to_check_it_0_cnu_36_in_5, msg_to_check_it_0_cnu_37_in_0, msg_to_check_it_0_cnu_37_in_1, msg_to_check_it_0_cnu_37_in_2, msg_to_check_it_0_cnu_37_in_3, msg_to_check_it_0_cnu_37_in_4, msg_to_check_it_0_cnu_37_in_5, msg_to_check_it_0_cnu_38_in_0, msg_to_check_it_0_cnu_38_in_1, msg_to_check_it_0_cnu_38_in_2, msg_to_check_it_0_cnu_38_in_3, msg_to_check_it_0_cnu_38_in_4, msg_to_check_it_0_cnu_38_in_5, msg_to_check_it_0_cnu_39_in_0, msg_to_check_it_0_cnu_39_in_1, msg_to_check_it_0_cnu_39_in_2, msg_to_check_it_0_cnu_39_in_3, msg_to_check_it_0_cnu_39_in_4, msg_to_check_it_0_cnu_39_in_5, msg_to_check_it_0_cnu_40_in_0, msg_to_check_it_0_cnu_40_in_1, msg_to_check_it_0_cnu_40_in_2, msg_to_check_it_0_cnu_40_in_3, msg_to_check_it_0_cnu_40_in_4, msg_to_check_it_0_cnu_40_in_5, msg_to_check_it_0_cnu_41_in_0, msg_to_check_it_0_cnu_41_in_1, msg_to_check_it_0_cnu_41_in_2, msg_to_check_it_0_cnu_41_in_3, msg_to_check_it_0_cnu_41_in_4, msg_to_check_it_0_cnu_41_in_5, msg_to_check_it_0_cnu_42_in_0, msg_to_check_it_0_cnu_42_in_1, msg_to_check_it_0_cnu_42_in_2, msg_to_check_it_0_cnu_42_in_3, msg_to_check_it_0_cnu_42_in_4, msg_to_check_it_0_cnu_42_in_5, msg_to_check_it_0_cnu_43_in_0, msg_to_check_it_0_cnu_43_in_1, msg_to_check_it_0_cnu_43_in_2, msg_to_check_it_0_cnu_43_in_3, msg_to_check_it_0_cnu_43_in_4, msg_to_check_it_0_cnu_43_in_5, msg_to_check_it_0_cnu_44_in_0, msg_to_check_it_0_cnu_44_in_1, msg_to_check_it_0_cnu_44_in_2, msg_to_check_it_0_cnu_44_in_3, msg_to_check_it_0_cnu_44_in_4, msg_to_check_it_0_cnu_44_in_5, msg_to_check_it_0_cnu_45_in_0, msg_to_check_it_0_cnu_45_in_1, msg_to_check_it_0_cnu_45_in_2, msg_to_check_it_0_cnu_45_in_3, msg_to_check_it_0_cnu_45_in_4, msg_to_check_it_0_cnu_45_in_5, msg_to_check_it_0_cnu_46_in_0, msg_to_check_it_0_cnu_46_in_1, msg_to_check_it_0_cnu_46_in_2, msg_to_check_it_0_cnu_46_in_3, msg_to_check_it_0_cnu_46_in_4, msg_to_check_it_0_cnu_46_in_5, msg_to_check_it_0_cnu_47_in_0, msg_to_check_it_0_cnu_47_in_1, msg_to_check_it_0_cnu_47_in_2, msg_to_check_it_0_cnu_47_in_3, msg_to_check_it_0_cnu_47_in_4, msg_to_check_it_0_cnu_47_in_5, msg_to_check_it_0_cnu_48_in_0, msg_to_check_it_0_cnu_48_in_1, msg_to_check_it_0_cnu_48_in_2, msg_to_check_it_0_cnu_48_in_3, msg_to_check_it_0_cnu_48_in_4, msg_to_check_it_0_cnu_48_in_5, msg_to_check_it_0_cnu_49_in_0, msg_to_check_it_0_cnu_49_in_1, msg_to_check_it_0_cnu_49_in_2, msg_to_check_it_0_cnu_49_in_3, msg_to_check_it_0_cnu_49_in_4, msg_to_check_it_0_cnu_49_in_5, msg_to_check_it_0_cnu_50_in_0, msg_to_check_it_0_cnu_50_in_1, msg_to_check_it_0_cnu_50_in_2, msg_to_check_it_0_cnu_50_in_3, msg_to_check_it_0_cnu_50_in_4, msg_to_check_it_0_cnu_50_in_5, msg_to_check_it_0_cnu_51_in_0, msg_to_check_it_0_cnu_51_in_1, msg_to_check_it_0_cnu_51_in_2, msg_to_check_it_0_cnu_51_in_3, msg_to_check_it_0_cnu_51_in_4, msg_to_check_it_0_cnu_51_in_5, msg_to_check_it_0_cnu_52_in_0, msg_to_check_it_0_cnu_52_in_1, msg_to_check_it_0_cnu_52_in_2, msg_to_check_it_0_cnu_52_in_3, msg_to_check_it_0_cnu_52_in_4, msg_to_check_it_0_cnu_52_in_5, msg_to_check_it_0_cnu_53_in_0, msg_to_check_it_0_cnu_53_in_1, msg_to_check_it_0_cnu_53_in_2, msg_to_check_it_0_cnu_53_in_3, msg_to_check_it_0_cnu_53_in_4, msg_to_check_it_0_cnu_53_in_5, msg_to_check_it_0_cnu_54_in_0, msg_to_check_it_0_cnu_54_in_1, msg_to_check_it_0_cnu_54_in_2, msg_to_check_it_0_cnu_54_in_3, msg_to_check_it_0_cnu_54_in_4, msg_to_check_it_0_cnu_54_in_5, msg_to_check_it_0_cnu_55_in_0, msg_to_check_it_0_cnu_55_in_1, msg_to_check_it_0_cnu_55_in_2, msg_to_check_it_0_cnu_55_in_3, msg_to_check_it_0_cnu_55_in_4, msg_to_check_it_0_cnu_55_in_5, msg_to_check_it_0_cnu_56_in_0, msg_to_check_it_0_cnu_56_in_1, msg_to_check_it_0_cnu_56_in_2, msg_to_check_it_0_cnu_56_in_3, msg_to_check_it_0_cnu_56_in_4, msg_to_check_it_0_cnu_56_in_5, msg_to_check_it_0_cnu_57_in_0, msg_to_check_it_0_cnu_57_in_1, msg_to_check_it_0_cnu_57_in_2, msg_to_check_it_0_cnu_57_in_3, msg_to_check_it_0_cnu_57_in_4, msg_to_check_it_0_cnu_57_in_5, msg_to_check_it_0_cnu_58_in_0, msg_to_check_it_0_cnu_58_in_1, msg_to_check_it_0_cnu_58_in_2, msg_to_check_it_0_cnu_58_in_3, msg_to_check_it_0_cnu_58_in_4, msg_to_check_it_0_cnu_58_in_5, msg_to_check_it_0_cnu_59_in_0, msg_to_check_it_0_cnu_59_in_1, msg_to_check_it_0_cnu_59_in_2, msg_to_check_it_0_cnu_59_in_3, msg_to_check_it_0_cnu_59_in_4, msg_to_check_it_0_cnu_59_in_5, msg_to_check_it_0_cnu_60_in_0, msg_to_check_it_0_cnu_60_in_1, msg_to_check_it_0_cnu_60_in_2, msg_to_check_it_0_cnu_60_in_3, msg_to_check_it_0_cnu_60_in_4, msg_to_check_it_0_cnu_60_in_5, msg_to_check_it_0_cnu_61_in_0, msg_to_check_it_0_cnu_61_in_1, msg_to_check_it_0_cnu_61_in_2, msg_to_check_it_0_cnu_61_in_3, msg_to_check_it_0_cnu_61_in_4, msg_to_check_it_0_cnu_61_in_5, msg_to_check_it_0_cnu_62_in_0, msg_to_check_it_0_cnu_62_in_1, msg_to_check_it_0_cnu_62_in_2, msg_to_check_it_0_cnu_62_in_3, msg_to_check_it_0_cnu_62_in_4, msg_to_check_it_0_cnu_62_in_5, msg_to_check_it_0_cnu_63_in_0, msg_to_check_it_0_cnu_63_in_1, msg_to_check_it_0_cnu_63_in_2, msg_to_check_it_0_cnu_63_in_3, msg_to_check_it_0_cnu_63_in_4, msg_to_check_it_0_cnu_63_in_5, msg_to_check_it_0_cnu_64_in_0, msg_to_check_it_0_cnu_64_in_1, msg_to_check_it_0_cnu_64_in_2, msg_to_check_it_0_cnu_64_in_3, msg_to_check_it_0_cnu_64_in_4, msg_to_check_it_0_cnu_64_in_5, msg_to_check_it_0_cnu_65_in_0, msg_to_check_it_0_cnu_65_in_1, msg_to_check_it_0_cnu_65_in_2, msg_to_check_it_0_cnu_65_in_3, msg_to_check_it_0_cnu_65_in_4, msg_to_check_it_0_cnu_65_in_5, msg_to_check_it_0_cnu_66_in_0, msg_to_check_it_0_cnu_66_in_1, msg_to_check_it_0_cnu_66_in_2, msg_to_check_it_0_cnu_66_in_3, msg_to_check_it_0_cnu_66_in_4, msg_to_check_it_0_cnu_66_in_5, msg_to_check_it_0_cnu_67_in_0, msg_to_check_it_0_cnu_67_in_1, msg_to_check_it_0_cnu_67_in_2, msg_to_check_it_0_cnu_67_in_3, msg_to_check_it_0_cnu_67_in_4, msg_to_check_it_0_cnu_67_in_5, msg_to_check_it_0_cnu_68_in_0, msg_to_check_it_0_cnu_68_in_1, msg_to_check_it_0_cnu_68_in_2, msg_to_check_it_0_cnu_68_in_3, msg_to_check_it_0_cnu_68_in_4, msg_to_check_it_0_cnu_68_in_5, msg_to_check_it_0_cnu_69_in_0, msg_to_check_it_0_cnu_69_in_1, msg_to_check_it_0_cnu_69_in_2, msg_to_check_it_0_cnu_69_in_3, msg_to_check_it_0_cnu_69_in_4, msg_to_check_it_0_cnu_69_in_5, msg_to_check_it_0_cnu_70_in_0, msg_to_check_it_0_cnu_70_in_1, msg_to_check_it_0_cnu_70_in_2, msg_to_check_it_0_cnu_70_in_3, msg_to_check_it_0_cnu_70_in_4, msg_to_check_it_0_cnu_70_in_5, msg_to_check_it_0_cnu_71_in_0, msg_to_check_it_0_cnu_71_in_1, msg_to_check_it_0_cnu_71_in_2, msg_to_check_it_0_cnu_71_in_3, msg_to_check_it_0_cnu_71_in_4, msg_to_check_it_0_cnu_71_in_5, msg_to_check_it_0_cnu_72_in_0, msg_to_check_it_0_cnu_72_in_1, msg_to_check_it_0_cnu_72_in_2, msg_to_check_it_0_cnu_72_in_3, msg_to_check_it_0_cnu_72_in_4, msg_to_check_it_0_cnu_72_in_5, msg_to_check_it_0_cnu_73_in_0, msg_to_check_it_0_cnu_73_in_1, msg_to_check_it_0_cnu_73_in_2, msg_to_check_it_0_cnu_73_in_3, msg_to_check_it_0_cnu_73_in_4, msg_to_check_it_0_cnu_73_in_5, msg_to_check_it_0_cnu_74_in_0, msg_to_check_it_0_cnu_74_in_1, msg_to_check_it_0_cnu_74_in_2, msg_to_check_it_0_cnu_74_in_3, msg_to_check_it_0_cnu_74_in_4, msg_to_check_it_0_cnu_74_in_5, msg_to_check_it_0_cnu_75_in_0, msg_to_check_it_0_cnu_75_in_1, msg_to_check_it_0_cnu_75_in_2, msg_to_check_it_0_cnu_75_in_3, msg_to_check_it_0_cnu_75_in_4, msg_to_check_it_0_cnu_75_in_5, msg_to_check_it_0_cnu_76_in_0, msg_to_check_it_0_cnu_76_in_1, msg_to_check_it_0_cnu_76_in_2, msg_to_check_it_0_cnu_76_in_3, msg_to_check_it_0_cnu_76_in_4, msg_to_check_it_0_cnu_76_in_5, msg_to_check_it_0_cnu_77_in_0, msg_to_check_it_0_cnu_77_in_1, msg_to_check_it_0_cnu_77_in_2, msg_to_check_it_0_cnu_77_in_3, msg_to_check_it_0_cnu_77_in_4, msg_to_check_it_0_cnu_77_in_5, msg_to_check_it_0_cnu_78_in_0, msg_to_check_it_0_cnu_78_in_1, msg_to_check_it_0_cnu_78_in_2, msg_to_check_it_0_cnu_78_in_3, msg_to_check_it_0_cnu_78_in_4, msg_to_check_it_0_cnu_78_in_5, msg_to_check_it_0_cnu_79_in_0, msg_to_check_it_0_cnu_79_in_1, msg_to_check_it_0_cnu_79_in_2, msg_to_check_it_0_cnu_79_in_3, msg_to_check_it_0_cnu_79_in_4, msg_to_check_it_0_cnu_79_in_5, msg_to_check_it_0_cnu_80_in_0, msg_to_check_it_0_cnu_80_in_1, msg_to_check_it_0_cnu_80_in_2, msg_to_check_it_0_cnu_80_in_3, msg_to_check_it_0_cnu_80_in_4, msg_to_check_it_0_cnu_80_in_5, msg_to_check_it_0_cnu_81_in_0, msg_to_check_it_0_cnu_81_in_1, msg_to_check_it_0_cnu_81_in_2, msg_to_check_it_0_cnu_81_in_3, msg_to_check_it_0_cnu_81_in_4, msg_to_check_it_0_cnu_81_in_5, msg_to_check_it_0_cnu_82_in_0, msg_to_check_it_0_cnu_82_in_1, msg_to_check_it_0_cnu_82_in_2, msg_to_check_it_0_cnu_82_in_3, msg_to_check_it_0_cnu_82_in_4, msg_to_check_it_0_cnu_82_in_5, msg_to_check_it_0_cnu_83_in_0, msg_to_check_it_0_cnu_83_in_1, msg_to_check_it_0_cnu_83_in_2, msg_to_check_it_0_cnu_83_in_3, msg_to_check_it_0_cnu_83_in_4, msg_to_check_it_0_cnu_83_in_5, msg_to_check_it_0_cnu_84_in_0, msg_to_check_it_0_cnu_84_in_1, msg_to_check_it_0_cnu_84_in_2, msg_to_check_it_0_cnu_84_in_3, msg_to_check_it_0_cnu_84_in_4, msg_to_check_it_0_cnu_84_in_5, msg_to_check_it_0_cnu_85_in_0, msg_to_check_it_0_cnu_85_in_1, msg_to_check_it_0_cnu_85_in_2, msg_to_check_it_0_cnu_85_in_3, msg_to_check_it_0_cnu_85_in_4, msg_to_check_it_0_cnu_85_in_5, msg_to_check_it_0_cnu_86_in_0, msg_to_check_it_0_cnu_86_in_1, msg_to_check_it_0_cnu_86_in_2, msg_to_check_it_0_cnu_86_in_3, msg_to_check_it_0_cnu_86_in_4, msg_to_check_it_0_cnu_86_in_5, msg_to_check_it_0_cnu_87_in_0, msg_to_check_it_0_cnu_87_in_1, msg_to_check_it_0_cnu_87_in_2, msg_to_check_it_0_cnu_87_in_3, msg_to_check_it_0_cnu_87_in_4, msg_to_check_it_0_cnu_87_in_5, msg_to_check_it_0_cnu_88_in_0, msg_to_check_it_0_cnu_88_in_1, msg_to_check_it_0_cnu_88_in_2, msg_to_check_it_0_cnu_88_in_3, msg_to_check_it_0_cnu_88_in_4, msg_to_check_it_0_cnu_88_in_5, msg_to_check_it_0_cnu_89_in_0, msg_to_check_it_0_cnu_89_in_1, msg_to_check_it_0_cnu_89_in_2, msg_to_check_it_0_cnu_89_in_3, msg_to_check_it_0_cnu_89_in_4, msg_to_check_it_0_cnu_89_in_5, msg_to_check_it_0_cnu_90_in_0, msg_to_check_it_0_cnu_90_in_1, msg_to_check_it_0_cnu_90_in_2, msg_to_check_it_0_cnu_90_in_3, msg_to_check_it_0_cnu_90_in_4, msg_to_check_it_0_cnu_90_in_5, msg_to_check_it_0_cnu_91_in_0, msg_to_check_it_0_cnu_91_in_1, msg_to_check_it_0_cnu_91_in_2, msg_to_check_it_0_cnu_91_in_3, msg_to_check_it_0_cnu_91_in_4, msg_to_check_it_0_cnu_91_in_5, msg_to_check_it_0_cnu_92_in_0, msg_to_check_it_0_cnu_92_in_1, msg_to_check_it_0_cnu_92_in_2, msg_to_check_it_0_cnu_92_in_3, msg_to_check_it_0_cnu_92_in_4, msg_to_check_it_0_cnu_92_in_5, msg_to_check_it_0_cnu_93_in_0, msg_to_check_it_0_cnu_93_in_1, msg_to_check_it_0_cnu_93_in_2, msg_to_check_it_0_cnu_93_in_3, msg_to_check_it_0_cnu_93_in_4, msg_to_check_it_0_cnu_93_in_5, msg_to_check_it_0_cnu_94_in_0, msg_to_check_it_0_cnu_94_in_1, msg_to_check_it_0_cnu_94_in_2, msg_to_check_it_0_cnu_94_in_3, msg_to_check_it_0_cnu_94_in_4, msg_to_check_it_0_cnu_94_in_5, msg_to_check_it_0_cnu_95_in_0, msg_to_check_it_0_cnu_95_in_1, msg_to_check_it_0_cnu_95_in_2, msg_to_check_it_0_cnu_95_in_3, msg_to_check_it_0_cnu_95_in_4, msg_to_check_it_0_cnu_95_in_5, msg_to_check_it_0_cnu_96_in_0, msg_to_check_it_0_cnu_96_in_1, msg_to_check_it_0_cnu_96_in_2, msg_to_check_it_0_cnu_96_in_3, msg_to_check_it_0_cnu_96_in_4, msg_to_check_it_0_cnu_96_in_5, msg_to_check_it_0_cnu_97_in_0, msg_to_check_it_0_cnu_97_in_1, msg_to_check_it_0_cnu_97_in_2, msg_to_check_it_0_cnu_97_in_3, msg_to_check_it_0_cnu_97_in_4, msg_to_check_it_0_cnu_97_in_5, msg_to_check_it_0_cnu_98_in_0, msg_to_check_it_0_cnu_98_in_1, msg_to_check_it_0_cnu_98_in_2, msg_to_check_it_0_cnu_98_in_3, msg_to_check_it_0_cnu_98_in_4, msg_to_check_it_0_cnu_98_in_5, msg_to_check_it_1_cnu_0_in_0, msg_to_check_it_1_cnu_0_in_1, msg_to_check_it_1_cnu_0_in_2, msg_to_check_it_1_cnu_0_in_3, msg_to_check_it_1_cnu_0_in_4, msg_to_check_it_1_cnu_0_in_5, msg_to_check_it_1_cnu_1_in_0, msg_to_check_it_1_cnu_1_in_1, msg_to_check_it_1_cnu_1_in_2, msg_to_check_it_1_cnu_1_in_3, msg_to_check_it_1_cnu_1_in_4, msg_to_check_it_1_cnu_1_in_5, msg_to_check_it_1_cnu_2_in_0, msg_to_check_it_1_cnu_2_in_1, msg_to_check_it_1_cnu_2_in_2, msg_to_check_it_1_cnu_2_in_3, msg_to_check_it_1_cnu_2_in_4, msg_to_check_it_1_cnu_2_in_5, msg_to_check_it_1_cnu_3_in_0, msg_to_check_it_1_cnu_3_in_1, msg_to_check_it_1_cnu_3_in_2, msg_to_check_it_1_cnu_3_in_3, msg_to_check_it_1_cnu_3_in_4, msg_to_check_it_1_cnu_3_in_5, msg_to_check_it_1_cnu_4_in_0, msg_to_check_it_1_cnu_4_in_1, msg_to_check_it_1_cnu_4_in_2, msg_to_check_it_1_cnu_4_in_3, msg_to_check_it_1_cnu_4_in_4, msg_to_check_it_1_cnu_4_in_5, msg_to_check_it_1_cnu_5_in_0, msg_to_check_it_1_cnu_5_in_1, msg_to_check_it_1_cnu_5_in_2, msg_to_check_it_1_cnu_5_in_3, msg_to_check_it_1_cnu_5_in_4, msg_to_check_it_1_cnu_5_in_5, msg_to_check_it_1_cnu_6_in_0, msg_to_check_it_1_cnu_6_in_1, msg_to_check_it_1_cnu_6_in_2, msg_to_check_it_1_cnu_6_in_3, msg_to_check_it_1_cnu_6_in_4, msg_to_check_it_1_cnu_6_in_5, msg_to_check_it_1_cnu_7_in_0, msg_to_check_it_1_cnu_7_in_1, msg_to_check_it_1_cnu_7_in_2, msg_to_check_it_1_cnu_7_in_3, msg_to_check_it_1_cnu_7_in_4, msg_to_check_it_1_cnu_7_in_5, msg_to_check_it_1_cnu_8_in_0, msg_to_check_it_1_cnu_8_in_1, msg_to_check_it_1_cnu_8_in_2, msg_to_check_it_1_cnu_8_in_3, msg_to_check_it_1_cnu_8_in_4, msg_to_check_it_1_cnu_8_in_5, msg_to_check_it_1_cnu_9_in_0, msg_to_check_it_1_cnu_9_in_1, msg_to_check_it_1_cnu_9_in_2, msg_to_check_it_1_cnu_9_in_3, msg_to_check_it_1_cnu_9_in_4, msg_to_check_it_1_cnu_9_in_5, msg_to_check_it_1_cnu_10_in_0, msg_to_check_it_1_cnu_10_in_1, msg_to_check_it_1_cnu_10_in_2, msg_to_check_it_1_cnu_10_in_3, msg_to_check_it_1_cnu_10_in_4, msg_to_check_it_1_cnu_10_in_5, msg_to_check_it_1_cnu_11_in_0, msg_to_check_it_1_cnu_11_in_1, msg_to_check_it_1_cnu_11_in_2, msg_to_check_it_1_cnu_11_in_3, msg_to_check_it_1_cnu_11_in_4, msg_to_check_it_1_cnu_11_in_5, msg_to_check_it_1_cnu_12_in_0, msg_to_check_it_1_cnu_12_in_1, msg_to_check_it_1_cnu_12_in_2, msg_to_check_it_1_cnu_12_in_3, msg_to_check_it_1_cnu_12_in_4, msg_to_check_it_1_cnu_12_in_5, msg_to_check_it_1_cnu_13_in_0, msg_to_check_it_1_cnu_13_in_1, msg_to_check_it_1_cnu_13_in_2, msg_to_check_it_1_cnu_13_in_3, msg_to_check_it_1_cnu_13_in_4, msg_to_check_it_1_cnu_13_in_5, msg_to_check_it_1_cnu_14_in_0, msg_to_check_it_1_cnu_14_in_1, msg_to_check_it_1_cnu_14_in_2, msg_to_check_it_1_cnu_14_in_3, msg_to_check_it_1_cnu_14_in_4, msg_to_check_it_1_cnu_14_in_5, msg_to_check_it_1_cnu_15_in_0, msg_to_check_it_1_cnu_15_in_1, msg_to_check_it_1_cnu_15_in_2, msg_to_check_it_1_cnu_15_in_3, msg_to_check_it_1_cnu_15_in_4, msg_to_check_it_1_cnu_15_in_5, msg_to_check_it_1_cnu_16_in_0, msg_to_check_it_1_cnu_16_in_1, msg_to_check_it_1_cnu_16_in_2, msg_to_check_it_1_cnu_16_in_3, msg_to_check_it_1_cnu_16_in_4, msg_to_check_it_1_cnu_16_in_5, msg_to_check_it_1_cnu_17_in_0, msg_to_check_it_1_cnu_17_in_1, msg_to_check_it_1_cnu_17_in_2, msg_to_check_it_1_cnu_17_in_3, msg_to_check_it_1_cnu_17_in_4, msg_to_check_it_1_cnu_17_in_5, msg_to_check_it_1_cnu_18_in_0, msg_to_check_it_1_cnu_18_in_1, msg_to_check_it_1_cnu_18_in_2, msg_to_check_it_1_cnu_18_in_3, msg_to_check_it_1_cnu_18_in_4, msg_to_check_it_1_cnu_18_in_5, msg_to_check_it_1_cnu_19_in_0, msg_to_check_it_1_cnu_19_in_1, msg_to_check_it_1_cnu_19_in_2, msg_to_check_it_1_cnu_19_in_3, msg_to_check_it_1_cnu_19_in_4, msg_to_check_it_1_cnu_19_in_5, msg_to_check_it_1_cnu_20_in_0, msg_to_check_it_1_cnu_20_in_1, msg_to_check_it_1_cnu_20_in_2, msg_to_check_it_1_cnu_20_in_3, msg_to_check_it_1_cnu_20_in_4, msg_to_check_it_1_cnu_20_in_5, msg_to_check_it_1_cnu_21_in_0, msg_to_check_it_1_cnu_21_in_1, msg_to_check_it_1_cnu_21_in_2, msg_to_check_it_1_cnu_21_in_3, msg_to_check_it_1_cnu_21_in_4, msg_to_check_it_1_cnu_21_in_5, msg_to_check_it_1_cnu_22_in_0, msg_to_check_it_1_cnu_22_in_1, msg_to_check_it_1_cnu_22_in_2, msg_to_check_it_1_cnu_22_in_3, msg_to_check_it_1_cnu_22_in_4, msg_to_check_it_1_cnu_22_in_5, msg_to_check_it_1_cnu_23_in_0, msg_to_check_it_1_cnu_23_in_1, msg_to_check_it_1_cnu_23_in_2, msg_to_check_it_1_cnu_23_in_3, msg_to_check_it_1_cnu_23_in_4, msg_to_check_it_1_cnu_23_in_5, msg_to_check_it_1_cnu_24_in_0, msg_to_check_it_1_cnu_24_in_1, msg_to_check_it_1_cnu_24_in_2, msg_to_check_it_1_cnu_24_in_3, msg_to_check_it_1_cnu_24_in_4, msg_to_check_it_1_cnu_24_in_5, msg_to_check_it_1_cnu_25_in_0, msg_to_check_it_1_cnu_25_in_1, msg_to_check_it_1_cnu_25_in_2, msg_to_check_it_1_cnu_25_in_3, msg_to_check_it_1_cnu_25_in_4, msg_to_check_it_1_cnu_25_in_5, msg_to_check_it_1_cnu_26_in_0, msg_to_check_it_1_cnu_26_in_1, msg_to_check_it_1_cnu_26_in_2, msg_to_check_it_1_cnu_26_in_3, msg_to_check_it_1_cnu_26_in_4, msg_to_check_it_1_cnu_26_in_5, msg_to_check_it_1_cnu_27_in_0, msg_to_check_it_1_cnu_27_in_1, msg_to_check_it_1_cnu_27_in_2, msg_to_check_it_1_cnu_27_in_3, msg_to_check_it_1_cnu_27_in_4, msg_to_check_it_1_cnu_27_in_5, msg_to_check_it_1_cnu_28_in_0, msg_to_check_it_1_cnu_28_in_1, msg_to_check_it_1_cnu_28_in_2, msg_to_check_it_1_cnu_28_in_3, msg_to_check_it_1_cnu_28_in_4, msg_to_check_it_1_cnu_28_in_5, msg_to_check_it_1_cnu_29_in_0, msg_to_check_it_1_cnu_29_in_1, msg_to_check_it_1_cnu_29_in_2, msg_to_check_it_1_cnu_29_in_3, msg_to_check_it_1_cnu_29_in_4, msg_to_check_it_1_cnu_29_in_5, msg_to_check_it_1_cnu_30_in_0, msg_to_check_it_1_cnu_30_in_1, msg_to_check_it_1_cnu_30_in_2, msg_to_check_it_1_cnu_30_in_3, msg_to_check_it_1_cnu_30_in_4, msg_to_check_it_1_cnu_30_in_5, msg_to_check_it_1_cnu_31_in_0, msg_to_check_it_1_cnu_31_in_1, msg_to_check_it_1_cnu_31_in_2, msg_to_check_it_1_cnu_31_in_3, msg_to_check_it_1_cnu_31_in_4, msg_to_check_it_1_cnu_31_in_5, msg_to_check_it_1_cnu_32_in_0, msg_to_check_it_1_cnu_32_in_1, msg_to_check_it_1_cnu_32_in_2, msg_to_check_it_1_cnu_32_in_3, msg_to_check_it_1_cnu_32_in_4, msg_to_check_it_1_cnu_32_in_5, msg_to_check_it_1_cnu_33_in_0, msg_to_check_it_1_cnu_33_in_1, msg_to_check_it_1_cnu_33_in_2, msg_to_check_it_1_cnu_33_in_3, msg_to_check_it_1_cnu_33_in_4, msg_to_check_it_1_cnu_33_in_5, msg_to_check_it_1_cnu_34_in_0, msg_to_check_it_1_cnu_34_in_1, msg_to_check_it_1_cnu_34_in_2, msg_to_check_it_1_cnu_34_in_3, msg_to_check_it_1_cnu_34_in_4, msg_to_check_it_1_cnu_34_in_5, msg_to_check_it_1_cnu_35_in_0, msg_to_check_it_1_cnu_35_in_1, msg_to_check_it_1_cnu_35_in_2, msg_to_check_it_1_cnu_35_in_3, msg_to_check_it_1_cnu_35_in_4, msg_to_check_it_1_cnu_35_in_5, msg_to_check_it_1_cnu_36_in_0, msg_to_check_it_1_cnu_36_in_1, msg_to_check_it_1_cnu_36_in_2, msg_to_check_it_1_cnu_36_in_3, msg_to_check_it_1_cnu_36_in_4, msg_to_check_it_1_cnu_36_in_5, msg_to_check_it_1_cnu_37_in_0, msg_to_check_it_1_cnu_37_in_1, msg_to_check_it_1_cnu_37_in_2, msg_to_check_it_1_cnu_37_in_3, msg_to_check_it_1_cnu_37_in_4, msg_to_check_it_1_cnu_37_in_5, msg_to_check_it_1_cnu_38_in_0, msg_to_check_it_1_cnu_38_in_1, msg_to_check_it_1_cnu_38_in_2, msg_to_check_it_1_cnu_38_in_3, msg_to_check_it_1_cnu_38_in_4, msg_to_check_it_1_cnu_38_in_5, msg_to_check_it_1_cnu_39_in_0, msg_to_check_it_1_cnu_39_in_1, msg_to_check_it_1_cnu_39_in_2, msg_to_check_it_1_cnu_39_in_3, msg_to_check_it_1_cnu_39_in_4, msg_to_check_it_1_cnu_39_in_5, msg_to_check_it_1_cnu_40_in_0, msg_to_check_it_1_cnu_40_in_1, msg_to_check_it_1_cnu_40_in_2, msg_to_check_it_1_cnu_40_in_3, msg_to_check_it_1_cnu_40_in_4, msg_to_check_it_1_cnu_40_in_5, msg_to_check_it_1_cnu_41_in_0, msg_to_check_it_1_cnu_41_in_1, msg_to_check_it_1_cnu_41_in_2, msg_to_check_it_1_cnu_41_in_3, msg_to_check_it_1_cnu_41_in_4, msg_to_check_it_1_cnu_41_in_5, msg_to_check_it_1_cnu_42_in_0, msg_to_check_it_1_cnu_42_in_1, msg_to_check_it_1_cnu_42_in_2, msg_to_check_it_1_cnu_42_in_3, msg_to_check_it_1_cnu_42_in_4, msg_to_check_it_1_cnu_42_in_5, msg_to_check_it_1_cnu_43_in_0, msg_to_check_it_1_cnu_43_in_1, msg_to_check_it_1_cnu_43_in_2, msg_to_check_it_1_cnu_43_in_3, msg_to_check_it_1_cnu_43_in_4, msg_to_check_it_1_cnu_43_in_5, msg_to_check_it_1_cnu_44_in_0, msg_to_check_it_1_cnu_44_in_1, msg_to_check_it_1_cnu_44_in_2, msg_to_check_it_1_cnu_44_in_3, msg_to_check_it_1_cnu_44_in_4, msg_to_check_it_1_cnu_44_in_5, msg_to_check_it_1_cnu_45_in_0, msg_to_check_it_1_cnu_45_in_1, msg_to_check_it_1_cnu_45_in_2, msg_to_check_it_1_cnu_45_in_3, msg_to_check_it_1_cnu_45_in_4, msg_to_check_it_1_cnu_45_in_5, msg_to_check_it_1_cnu_46_in_0, msg_to_check_it_1_cnu_46_in_1, msg_to_check_it_1_cnu_46_in_2, msg_to_check_it_1_cnu_46_in_3, msg_to_check_it_1_cnu_46_in_4, msg_to_check_it_1_cnu_46_in_5, msg_to_check_it_1_cnu_47_in_0, msg_to_check_it_1_cnu_47_in_1, msg_to_check_it_1_cnu_47_in_2, msg_to_check_it_1_cnu_47_in_3, msg_to_check_it_1_cnu_47_in_4, msg_to_check_it_1_cnu_47_in_5, msg_to_check_it_1_cnu_48_in_0, msg_to_check_it_1_cnu_48_in_1, msg_to_check_it_1_cnu_48_in_2, msg_to_check_it_1_cnu_48_in_3, msg_to_check_it_1_cnu_48_in_4, msg_to_check_it_1_cnu_48_in_5, msg_to_check_it_1_cnu_49_in_0, msg_to_check_it_1_cnu_49_in_1, msg_to_check_it_1_cnu_49_in_2, msg_to_check_it_1_cnu_49_in_3, msg_to_check_it_1_cnu_49_in_4, msg_to_check_it_1_cnu_49_in_5, msg_to_check_it_1_cnu_50_in_0, msg_to_check_it_1_cnu_50_in_1, msg_to_check_it_1_cnu_50_in_2, msg_to_check_it_1_cnu_50_in_3, msg_to_check_it_1_cnu_50_in_4, msg_to_check_it_1_cnu_50_in_5, msg_to_check_it_1_cnu_51_in_0, msg_to_check_it_1_cnu_51_in_1, msg_to_check_it_1_cnu_51_in_2, msg_to_check_it_1_cnu_51_in_3, msg_to_check_it_1_cnu_51_in_4, msg_to_check_it_1_cnu_51_in_5, msg_to_check_it_1_cnu_52_in_0, msg_to_check_it_1_cnu_52_in_1, msg_to_check_it_1_cnu_52_in_2, msg_to_check_it_1_cnu_52_in_3, msg_to_check_it_1_cnu_52_in_4, msg_to_check_it_1_cnu_52_in_5, msg_to_check_it_1_cnu_53_in_0, msg_to_check_it_1_cnu_53_in_1, msg_to_check_it_1_cnu_53_in_2, msg_to_check_it_1_cnu_53_in_3, msg_to_check_it_1_cnu_53_in_4, msg_to_check_it_1_cnu_53_in_5, msg_to_check_it_1_cnu_54_in_0, msg_to_check_it_1_cnu_54_in_1, msg_to_check_it_1_cnu_54_in_2, msg_to_check_it_1_cnu_54_in_3, msg_to_check_it_1_cnu_54_in_4, msg_to_check_it_1_cnu_54_in_5, msg_to_check_it_1_cnu_55_in_0, msg_to_check_it_1_cnu_55_in_1, msg_to_check_it_1_cnu_55_in_2, msg_to_check_it_1_cnu_55_in_3, msg_to_check_it_1_cnu_55_in_4, msg_to_check_it_1_cnu_55_in_5, msg_to_check_it_1_cnu_56_in_0, msg_to_check_it_1_cnu_56_in_1, msg_to_check_it_1_cnu_56_in_2, msg_to_check_it_1_cnu_56_in_3, msg_to_check_it_1_cnu_56_in_4, msg_to_check_it_1_cnu_56_in_5, msg_to_check_it_1_cnu_57_in_0, msg_to_check_it_1_cnu_57_in_1, msg_to_check_it_1_cnu_57_in_2, msg_to_check_it_1_cnu_57_in_3, msg_to_check_it_1_cnu_57_in_4, msg_to_check_it_1_cnu_57_in_5, msg_to_check_it_1_cnu_58_in_0, msg_to_check_it_1_cnu_58_in_1, msg_to_check_it_1_cnu_58_in_2, msg_to_check_it_1_cnu_58_in_3, msg_to_check_it_1_cnu_58_in_4, msg_to_check_it_1_cnu_58_in_5, msg_to_check_it_1_cnu_59_in_0, msg_to_check_it_1_cnu_59_in_1, msg_to_check_it_1_cnu_59_in_2, msg_to_check_it_1_cnu_59_in_3, msg_to_check_it_1_cnu_59_in_4, msg_to_check_it_1_cnu_59_in_5, msg_to_check_it_1_cnu_60_in_0, msg_to_check_it_1_cnu_60_in_1, msg_to_check_it_1_cnu_60_in_2, msg_to_check_it_1_cnu_60_in_3, msg_to_check_it_1_cnu_60_in_4, msg_to_check_it_1_cnu_60_in_5, msg_to_check_it_1_cnu_61_in_0, msg_to_check_it_1_cnu_61_in_1, msg_to_check_it_1_cnu_61_in_2, msg_to_check_it_1_cnu_61_in_3, msg_to_check_it_1_cnu_61_in_4, msg_to_check_it_1_cnu_61_in_5, msg_to_check_it_1_cnu_62_in_0, msg_to_check_it_1_cnu_62_in_1, msg_to_check_it_1_cnu_62_in_2, msg_to_check_it_1_cnu_62_in_3, msg_to_check_it_1_cnu_62_in_4, msg_to_check_it_1_cnu_62_in_5, msg_to_check_it_1_cnu_63_in_0, msg_to_check_it_1_cnu_63_in_1, msg_to_check_it_1_cnu_63_in_2, msg_to_check_it_1_cnu_63_in_3, msg_to_check_it_1_cnu_63_in_4, msg_to_check_it_1_cnu_63_in_5, msg_to_check_it_1_cnu_64_in_0, msg_to_check_it_1_cnu_64_in_1, msg_to_check_it_1_cnu_64_in_2, msg_to_check_it_1_cnu_64_in_3, msg_to_check_it_1_cnu_64_in_4, msg_to_check_it_1_cnu_64_in_5, msg_to_check_it_1_cnu_65_in_0, msg_to_check_it_1_cnu_65_in_1, msg_to_check_it_1_cnu_65_in_2, msg_to_check_it_1_cnu_65_in_3, msg_to_check_it_1_cnu_65_in_4, msg_to_check_it_1_cnu_65_in_5, msg_to_check_it_1_cnu_66_in_0, msg_to_check_it_1_cnu_66_in_1, msg_to_check_it_1_cnu_66_in_2, msg_to_check_it_1_cnu_66_in_3, msg_to_check_it_1_cnu_66_in_4, msg_to_check_it_1_cnu_66_in_5, msg_to_check_it_1_cnu_67_in_0, msg_to_check_it_1_cnu_67_in_1, msg_to_check_it_1_cnu_67_in_2, msg_to_check_it_1_cnu_67_in_3, msg_to_check_it_1_cnu_67_in_4, msg_to_check_it_1_cnu_67_in_5, msg_to_check_it_1_cnu_68_in_0, msg_to_check_it_1_cnu_68_in_1, msg_to_check_it_1_cnu_68_in_2, msg_to_check_it_1_cnu_68_in_3, msg_to_check_it_1_cnu_68_in_4, msg_to_check_it_1_cnu_68_in_5, msg_to_check_it_1_cnu_69_in_0, msg_to_check_it_1_cnu_69_in_1, msg_to_check_it_1_cnu_69_in_2, msg_to_check_it_1_cnu_69_in_3, msg_to_check_it_1_cnu_69_in_4, msg_to_check_it_1_cnu_69_in_5, msg_to_check_it_1_cnu_70_in_0, msg_to_check_it_1_cnu_70_in_1, msg_to_check_it_1_cnu_70_in_2, msg_to_check_it_1_cnu_70_in_3, msg_to_check_it_1_cnu_70_in_4, msg_to_check_it_1_cnu_70_in_5, msg_to_check_it_1_cnu_71_in_0, msg_to_check_it_1_cnu_71_in_1, msg_to_check_it_1_cnu_71_in_2, msg_to_check_it_1_cnu_71_in_3, msg_to_check_it_1_cnu_71_in_4, msg_to_check_it_1_cnu_71_in_5, msg_to_check_it_1_cnu_72_in_0, msg_to_check_it_1_cnu_72_in_1, msg_to_check_it_1_cnu_72_in_2, msg_to_check_it_1_cnu_72_in_3, msg_to_check_it_1_cnu_72_in_4, msg_to_check_it_1_cnu_72_in_5, msg_to_check_it_1_cnu_73_in_0, msg_to_check_it_1_cnu_73_in_1, msg_to_check_it_1_cnu_73_in_2, msg_to_check_it_1_cnu_73_in_3, msg_to_check_it_1_cnu_73_in_4, msg_to_check_it_1_cnu_73_in_5, msg_to_check_it_1_cnu_74_in_0, msg_to_check_it_1_cnu_74_in_1, msg_to_check_it_1_cnu_74_in_2, msg_to_check_it_1_cnu_74_in_3, msg_to_check_it_1_cnu_74_in_4, msg_to_check_it_1_cnu_74_in_5, msg_to_check_it_1_cnu_75_in_0, msg_to_check_it_1_cnu_75_in_1, msg_to_check_it_1_cnu_75_in_2, msg_to_check_it_1_cnu_75_in_3, msg_to_check_it_1_cnu_75_in_4, msg_to_check_it_1_cnu_75_in_5, msg_to_check_it_1_cnu_76_in_0, msg_to_check_it_1_cnu_76_in_1, msg_to_check_it_1_cnu_76_in_2, msg_to_check_it_1_cnu_76_in_3, msg_to_check_it_1_cnu_76_in_4, msg_to_check_it_1_cnu_76_in_5, msg_to_check_it_1_cnu_77_in_0, msg_to_check_it_1_cnu_77_in_1, msg_to_check_it_1_cnu_77_in_2, msg_to_check_it_1_cnu_77_in_3, msg_to_check_it_1_cnu_77_in_4, msg_to_check_it_1_cnu_77_in_5, msg_to_check_it_1_cnu_78_in_0, msg_to_check_it_1_cnu_78_in_1, msg_to_check_it_1_cnu_78_in_2, msg_to_check_it_1_cnu_78_in_3, msg_to_check_it_1_cnu_78_in_4, msg_to_check_it_1_cnu_78_in_5, msg_to_check_it_1_cnu_79_in_0, msg_to_check_it_1_cnu_79_in_1, msg_to_check_it_1_cnu_79_in_2, msg_to_check_it_1_cnu_79_in_3, msg_to_check_it_1_cnu_79_in_4, msg_to_check_it_1_cnu_79_in_5, msg_to_check_it_1_cnu_80_in_0, msg_to_check_it_1_cnu_80_in_1, msg_to_check_it_1_cnu_80_in_2, msg_to_check_it_1_cnu_80_in_3, msg_to_check_it_1_cnu_80_in_4, msg_to_check_it_1_cnu_80_in_5, msg_to_check_it_1_cnu_81_in_0, msg_to_check_it_1_cnu_81_in_1, msg_to_check_it_1_cnu_81_in_2, msg_to_check_it_1_cnu_81_in_3, msg_to_check_it_1_cnu_81_in_4, msg_to_check_it_1_cnu_81_in_5, msg_to_check_it_1_cnu_82_in_0, msg_to_check_it_1_cnu_82_in_1, msg_to_check_it_1_cnu_82_in_2, msg_to_check_it_1_cnu_82_in_3, msg_to_check_it_1_cnu_82_in_4, msg_to_check_it_1_cnu_82_in_5, msg_to_check_it_1_cnu_83_in_0, msg_to_check_it_1_cnu_83_in_1, msg_to_check_it_1_cnu_83_in_2, msg_to_check_it_1_cnu_83_in_3, msg_to_check_it_1_cnu_83_in_4, msg_to_check_it_1_cnu_83_in_5, msg_to_check_it_1_cnu_84_in_0, msg_to_check_it_1_cnu_84_in_1, msg_to_check_it_1_cnu_84_in_2, msg_to_check_it_1_cnu_84_in_3, msg_to_check_it_1_cnu_84_in_4, msg_to_check_it_1_cnu_84_in_5, msg_to_check_it_1_cnu_85_in_0, msg_to_check_it_1_cnu_85_in_1, msg_to_check_it_1_cnu_85_in_2, msg_to_check_it_1_cnu_85_in_3, msg_to_check_it_1_cnu_85_in_4, msg_to_check_it_1_cnu_85_in_5, msg_to_check_it_1_cnu_86_in_0, msg_to_check_it_1_cnu_86_in_1, msg_to_check_it_1_cnu_86_in_2, msg_to_check_it_1_cnu_86_in_3, msg_to_check_it_1_cnu_86_in_4, msg_to_check_it_1_cnu_86_in_5, msg_to_check_it_1_cnu_87_in_0, msg_to_check_it_1_cnu_87_in_1, msg_to_check_it_1_cnu_87_in_2, msg_to_check_it_1_cnu_87_in_3, msg_to_check_it_1_cnu_87_in_4, msg_to_check_it_1_cnu_87_in_5, msg_to_check_it_1_cnu_88_in_0, msg_to_check_it_1_cnu_88_in_1, msg_to_check_it_1_cnu_88_in_2, msg_to_check_it_1_cnu_88_in_3, msg_to_check_it_1_cnu_88_in_4, msg_to_check_it_1_cnu_88_in_5, msg_to_check_it_1_cnu_89_in_0, msg_to_check_it_1_cnu_89_in_1, msg_to_check_it_1_cnu_89_in_2, msg_to_check_it_1_cnu_89_in_3, msg_to_check_it_1_cnu_89_in_4, msg_to_check_it_1_cnu_89_in_5, msg_to_check_it_1_cnu_90_in_0, msg_to_check_it_1_cnu_90_in_1, msg_to_check_it_1_cnu_90_in_2, msg_to_check_it_1_cnu_90_in_3, msg_to_check_it_1_cnu_90_in_4, msg_to_check_it_1_cnu_90_in_5, msg_to_check_it_1_cnu_91_in_0, msg_to_check_it_1_cnu_91_in_1, msg_to_check_it_1_cnu_91_in_2, msg_to_check_it_1_cnu_91_in_3, msg_to_check_it_1_cnu_91_in_4, msg_to_check_it_1_cnu_91_in_5, msg_to_check_it_1_cnu_92_in_0, msg_to_check_it_1_cnu_92_in_1, msg_to_check_it_1_cnu_92_in_2, msg_to_check_it_1_cnu_92_in_3, msg_to_check_it_1_cnu_92_in_4, msg_to_check_it_1_cnu_92_in_5, msg_to_check_it_1_cnu_93_in_0, msg_to_check_it_1_cnu_93_in_1, msg_to_check_it_1_cnu_93_in_2, msg_to_check_it_1_cnu_93_in_3, msg_to_check_it_1_cnu_93_in_4, msg_to_check_it_1_cnu_93_in_5, msg_to_check_it_1_cnu_94_in_0, msg_to_check_it_1_cnu_94_in_1, msg_to_check_it_1_cnu_94_in_2, msg_to_check_it_1_cnu_94_in_3, msg_to_check_it_1_cnu_94_in_4, msg_to_check_it_1_cnu_94_in_5, msg_to_check_it_1_cnu_95_in_0, msg_to_check_it_1_cnu_95_in_1, msg_to_check_it_1_cnu_95_in_2, msg_to_check_it_1_cnu_95_in_3, msg_to_check_it_1_cnu_95_in_4, msg_to_check_it_1_cnu_95_in_5, msg_to_check_it_1_cnu_96_in_0, msg_to_check_it_1_cnu_96_in_1, msg_to_check_it_1_cnu_96_in_2, msg_to_check_it_1_cnu_96_in_3, msg_to_check_it_1_cnu_96_in_4, msg_to_check_it_1_cnu_96_in_5, msg_to_check_it_1_cnu_97_in_0, msg_to_check_it_1_cnu_97_in_1, msg_to_check_it_1_cnu_97_in_2, msg_to_check_it_1_cnu_97_in_3, msg_to_check_it_1_cnu_97_in_4, msg_to_check_it_1_cnu_97_in_5, msg_to_check_it_1_cnu_98_in_0, msg_to_check_it_1_cnu_98_in_1, msg_to_check_it_1_cnu_98_in_2, msg_to_check_it_1_cnu_98_in_3, msg_to_check_it_1_cnu_98_in_4, msg_to_check_it_1_cnu_98_in_5, msg_to_check_it_2_cnu_0_in_0, msg_to_check_it_2_cnu_0_in_1, msg_to_check_it_2_cnu_0_in_2, msg_to_check_it_2_cnu_0_in_3, msg_to_check_it_2_cnu_0_in_4, msg_to_check_it_2_cnu_0_in_5, msg_to_check_it_2_cnu_1_in_0, msg_to_check_it_2_cnu_1_in_1, msg_to_check_it_2_cnu_1_in_2, msg_to_check_it_2_cnu_1_in_3, msg_to_check_it_2_cnu_1_in_4, msg_to_check_it_2_cnu_1_in_5, msg_to_check_it_2_cnu_2_in_0, msg_to_check_it_2_cnu_2_in_1, msg_to_check_it_2_cnu_2_in_2, msg_to_check_it_2_cnu_2_in_3, msg_to_check_it_2_cnu_2_in_4, msg_to_check_it_2_cnu_2_in_5, msg_to_check_it_2_cnu_3_in_0, msg_to_check_it_2_cnu_3_in_1, msg_to_check_it_2_cnu_3_in_2, msg_to_check_it_2_cnu_3_in_3, msg_to_check_it_2_cnu_3_in_4, msg_to_check_it_2_cnu_3_in_5, msg_to_check_it_2_cnu_4_in_0, msg_to_check_it_2_cnu_4_in_1, msg_to_check_it_2_cnu_4_in_2, msg_to_check_it_2_cnu_4_in_3, msg_to_check_it_2_cnu_4_in_4, msg_to_check_it_2_cnu_4_in_5, msg_to_check_it_2_cnu_5_in_0, msg_to_check_it_2_cnu_5_in_1, msg_to_check_it_2_cnu_5_in_2, msg_to_check_it_2_cnu_5_in_3, msg_to_check_it_2_cnu_5_in_4, msg_to_check_it_2_cnu_5_in_5, msg_to_check_it_2_cnu_6_in_0, msg_to_check_it_2_cnu_6_in_1, msg_to_check_it_2_cnu_6_in_2, msg_to_check_it_2_cnu_6_in_3, msg_to_check_it_2_cnu_6_in_4, msg_to_check_it_2_cnu_6_in_5, msg_to_check_it_2_cnu_7_in_0, msg_to_check_it_2_cnu_7_in_1, msg_to_check_it_2_cnu_7_in_2, msg_to_check_it_2_cnu_7_in_3, msg_to_check_it_2_cnu_7_in_4, msg_to_check_it_2_cnu_7_in_5, msg_to_check_it_2_cnu_8_in_0, msg_to_check_it_2_cnu_8_in_1, msg_to_check_it_2_cnu_8_in_2, msg_to_check_it_2_cnu_8_in_3, msg_to_check_it_2_cnu_8_in_4, msg_to_check_it_2_cnu_8_in_5, msg_to_check_it_2_cnu_9_in_0, msg_to_check_it_2_cnu_9_in_1, msg_to_check_it_2_cnu_9_in_2, msg_to_check_it_2_cnu_9_in_3, msg_to_check_it_2_cnu_9_in_4, msg_to_check_it_2_cnu_9_in_5, msg_to_check_it_2_cnu_10_in_0, msg_to_check_it_2_cnu_10_in_1, msg_to_check_it_2_cnu_10_in_2, msg_to_check_it_2_cnu_10_in_3, msg_to_check_it_2_cnu_10_in_4, msg_to_check_it_2_cnu_10_in_5, msg_to_check_it_2_cnu_11_in_0, msg_to_check_it_2_cnu_11_in_1, msg_to_check_it_2_cnu_11_in_2, msg_to_check_it_2_cnu_11_in_3, msg_to_check_it_2_cnu_11_in_4, msg_to_check_it_2_cnu_11_in_5, msg_to_check_it_2_cnu_12_in_0, msg_to_check_it_2_cnu_12_in_1, msg_to_check_it_2_cnu_12_in_2, msg_to_check_it_2_cnu_12_in_3, msg_to_check_it_2_cnu_12_in_4, msg_to_check_it_2_cnu_12_in_5, msg_to_check_it_2_cnu_13_in_0, msg_to_check_it_2_cnu_13_in_1, msg_to_check_it_2_cnu_13_in_2, msg_to_check_it_2_cnu_13_in_3, msg_to_check_it_2_cnu_13_in_4, msg_to_check_it_2_cnu_13_in_5, msg_to_check_it_2_cnu_14_in_0, msg_to_check_it_2_cnu_14_in_1, msg_to_check_it_2_cnu_14_in_2, msg_to_check_it_2_cnu_14_in_3, msg_to_check_it_2_cnu_14_in_4, msg_to_check_it_2_cnu_14_in_5, msg_to_check_it_2_cnu_15_in_0, msg_to_check_it_2_cnu_15_in_1, msg_to_check_it_2_cnu_15_in_2, msg_to_check_it_2_cnu_15_in_3, msg_to_check_it_2_cnu_15_in_4, msg_to_check_it_2_cnu_15_in_5, msg_to_check_it_2_cnu_16_in_0, msg_to_check_it_2_cnu_16_in_1, msg_to_check_it_2_cnu_16_in_2, msg_to_check_it_2_cnu_16_in_3, msg_to_check_it_2_cnu_16_in_4, msg_to_check_it_2_cnu_16_in_5, msg_to_check_it_2_cnu_17_in_0, msg_to_check_it_2_cnu_17_in_1, msg_to_check_it_2_cnu_17_in_2, msg_to_check_it_2_cnu_17_in_3, msg_to_check_it_2_cnu_17_in_4, msg_to_check_it_2_cnu_17_in_5, msg_to_check_it_2_cnu_18_in_0, msg_to_check_it_2_cnu_18_in_1, msg_to_check_it_2_cnu_18_in_2, msg_to_check_it_2_cnu_18_in_3, msg_to_check_it_2_cnu_18_in_4, msg_to_check_it_2_cnu_18_in_5, msg_to_check_it_2_cnu_19_in_0, msg_to_check_it_2_cnu_19_in_1, msg_to_check_it_2_cnu_19_in_2, msg_to_check_it_2_cnu_19_in_3, msg_to_check_it_2_cnu_19_in_4, msg_to_check_it_2_cnu_19_in_5, msg_to_check_it_2_cnu_20_in_0, msg_to_check_it_2_cnu_20_in_1, msg_to_check_it_2_cnu_20_in_2, msg_to_check_it_2_cnu_20_in_3, msg_to_check_it_2_cnu_20_in_4, msg_to_check_it_2_cnu_20_in_5, msg_to_check_it_2_cnu_21_in_0, msg_to_check_it_2_cnu_21_in_1, msg_to_check_it_2_cnu_21_in_2, msg_to_check_it_2_cnu_21_in_3, msg_to_check_it_2_cnu_21_in_4, msg_to_check_it_2_cnu_21_in_5, msg_to_check_it_2_cnu_22_in_0, msg_to_check_it_2_cnu_22_in_1, msg_to_check_it_2_cnu_22_in_2, msg_to_check_it_2_cnu_22_in_3, msg_to_check_it_2_cnu_22_in_4, msg_to_check_it_2_cnu_22_in_5, msg_to_check_it_2_cnu_23_in_0, msg_to_check_it_2_cnu_23_in_1, msg_to_check_it_2_cnu_23_in_2, msg_to_check_it_2_cnu_23_in_3, msg_to_check_it_2_cnu_23_in_4, msg_to_check_it_2_cnu_23_in_5, msg_to_check_it_2_cnu_24_in_0, msg_to_check_it_2_cnu_24_in_1, msg_to_check_it_2_cnu_24_in_2, msg_to_check_it_2_cnu_24_in_3, msg_to_check_it_2_cnu_24_in_4, msg_to_check_it_2_cnu_24_in_5, msg_to_check_it_2_cnu_25_in_0, msg_to_check_it_2_cnu_25_in_1, msg_to_check_it_2_cnu_25_in_2, msg_to_check_it_2_cnu_25_in_3, msg_to_check_it_2_cnu_25_in_4, msg_to_check_it_2_cnu_25_in_5, msg_to_check_it_2_cnu_26_in_0, msg_to_check_it_2_cnu_26_in_1, msg_to_check_it_2_cnu_26_in_2, msg_to_check_it_2_cnu_26_in_3, msg_to_check_it_2_cnu_26_in_4, msg_to_check_it_2_cnu_26_in_5, msg_to_check_it_2_cnu_27_in_0, msg_to_check_it_2_cnu_27_in_1, msg_to_check_it_2_cnu_27_in_2, msg_to_check_it_2_cnu_27_in_3, msg_to_check_it_2_cnu_27_in_4, msg_to_check_it_2_cnu_27_in_5, msg_to_check_it_2_cnu_28_in_0, msg_to_check_it_2_cnu_28_in_1, msg_to_check_it_2_cnu_28_in_2, msg_to_check_it_2_cnu_28_in_3, msg_to_check_it_2_cnu_28_in_4, msg_to_check_it_2_cnu_28_in_5, msg_to_check_it_2_cnu_29_in_0, msg_to_check_it_2_cnu_29_in_1, msg_to_check_it_2_cnu_29_in_2, msg_to_check_it_2_cnu_29_in_3, msg_to_check_it_2_cnu_29_in_4, msg_to_check_it_2_cnu_29_in_5, msg_to_check_it_2_cnu_30_in_0, msg_to_check_it_2_cnu_30_in_1, msg_to_check_it_2_cnu_30_in_2, msg_to_check_it_2_cnu_30_in_3, msg_to_check_it_2_cnu_30_in_4, msg_to_check_it_2_cnu_30_in_5, msg_to_check_it_2_cnu_31_in_0, msg_to_check_it_2_cnu_31_in_1, msg_to_check_it_2_cnu_31_in_2, msg_to_check_it_2_cnu_31_in_3, msg_to_check_it_2_cnu_31_in_4, msg_to_check_it_2_cnu_31_in_5, msg_to_check_it_2_cnu_32_in_0, msg_to_check_it_2_cnu_32_in_1, msg_to_check_it_2_cnu_32_in_2, msg_to_check_it_2_cnu_32_in_3, msg_to_check_it_2_cnu_32_in_4, msg_to_check_it_2_cnu_32_in_5, msg_to_check_it_2_cnu_33_in_0, msg_to_check_it_2_cnu_33_in_1, msg_to_check_it_2_cnu_33_in_2, msg_to_check_it_2_cnu_33_in_3, msg_to_check_it_2_cnu_33_in_4, msg_to_check_it_2_cnu_33_in_5, msg_to_check_it_2_cnu_34_in_0, msg_to_check_it_2_cnu_34_in_1, msg_to_check_it_2_cnu_34_in_2, msg_to_check_it_2_cnu_34_in_3, msg_to_check_it_2_cnu_34_in_4, msg_to_check_it_2_cnu_34_in_5, msg_to_check_it_2_cnu_35_in_0, msg_to_check_it_2_cnu_35_in_1, msg_to_check_it_2_cnu_35_in_2, msg_to_check_it_2_cnu_35_in_3, msg_to_check_it_2_cnu_35_in_4, msg_to_check_it_2_cnu_35_in_5, msg_to_check_it_2_cnu_36_in_0, msg_to_check_it_2_cnu_36_in_1, msg_to_check_it_2_cnu_36_in_2, msg_to_check_it_2_cnu_36_in_3, msg_to_check_it_2_cnu_36_in_4, msg_to_check_it_2_cnu_36_in_5, msg_to_check_it_2_cnu_37_in_0, msg_to_check_it_2_cnu_37_in_1, msg_to_check_it_2_cnu_37_in_2, msg_to_check_it_2_cnu_37_in_3, msg_to_check_it_2_cnu_37_in_4, msg_to_check_it_2_cnu_37_in_5, msg_to_check_it_2_cnu_38_in_0, msg_to_check_it_2_cnu_38_in_1, msg_to_check_it_2_cnu_38_in_2, msg_to_check_it_2_cnu_38_in_3, msg_to_check_it_2_cnu_38_in_4, msg_to_check_it_2_cnu_38_in_5, msg_to_check_it_2_cnu_39_in_0, msg_to_check_it_2_cnu_39_in_1, msg_to_check_it_2_cnu_39_in_2, msg_to_check_it_2_cnu_39_in_3, msg_to_check_it_2_cnu_39_in_4, msg_to_check_it_2_cnu_39_in_5, msg_to_check_it_2_cnu_40_in_0, msg_to_check_it_2_cnu_40_in_1, msg_to_check_it_2_cnu_40_in_2, msg_to_check_it_2_cnu_40_in_3, msg_to_check_it_2_cnu_40_in_4, msg_to_check_it_2_cnu_40_in_5, msg_to_check_it_2_cnu_41_in_0, msg_to_check_it_2_cnu_41_in_1, msg_to_check_it_2_cnu_41_in_2, msg_to_check_it_2_cnu_41_in_3, msg_to_check_it_2_cnu_41_in_4, msg_to_check_it_2_cnu_41_in_5, msg_to_check_it_2_cnu_42_in_0, msg_to_check_it_2_cnu_42_in_1, msg_to_check_it_2_cnu_42_in_2, msg_to_check_it_2_cnu_42_in_3, msg_to_check_it_2_cnu_42_in_4, msg_to_check_it_2_cnu_42_in_5, msg_to_check_it_2_cnu_43_in_0, msg_to_check_it_2_cnu_43_in_1, msg_to_check_it_2_cnu_43_in_2, msg_to_check_it_2_cnu_43_in_3, msg_to_check_it_2_cnu_43_in_4, msg_to_check_it_2_cnu_43_in_5, msg_to_check_it_2_cnu_44_in_0, msg_to_check_it_2_cnu_44_in_1, msg_to_check_it_2_cnu_44_in_2, msg_to_check_it_2_cnu_44_in_3, msg_to_check_it_2_cnu_44_in_4, msg_to_check_it_2_cnu_44_in_5, msg_to_check_it_2_cnu_45_in_0, msg_to_check_it_2_cnu_45_in_1, msg_to_check_it_2_cnu_45_in_2, msg_to_check_it_2_cnu_45_in_3, msg_to_check_it_2_cnu_45_in_4, msg_to_check_it_2_cnu_45_in_5, msg_to_check_it_2_cnu_46_in_0, msg_to_check_it_2_cnu_46_in_1, msg_to_check_it_2_cnu_46_in_2, msg_to_check_it_2_cnu_46_in_3, msg_to_check_it_2_cnu_46_in_4, msg_to_check_it_2_cnu_46_in_5, msg_to_check_it_2_cnu_47_in_0, msg_to_check_it_2_cnu_47_in_1, msg_to_check_it_2_cnu_47_in_2, msg_to_check_it_2_cnu_47_in_3, msg_to_check_it_2_cnu_47_in_4, msg_to_check_it_2_cnu_47_in_5, msg_to_check_it_2_cnu_48_in_0, msg_to_check_it_2_cnu_48_in_1, msg_to_check_it_2_cnu_48_in_2, msg_to_check_it_2_cnu_48_in_3, msg_to_check_it_2_cnu_48_in_4, msg_to_check_it_2_cnu_48_in_5, msg_to_check_it_2_cnu_49_in_0, msg_to_check_it_2_cnu_49_in_1, msg_to_check_it_2_cnu_49_in_2, msg_to_check_it_2_cnu_49_in_3, msg_to_check_it_2_cnu_49_in_4, msg_to_check_it_2_cnu_49_in_5, msg_to_check_it_2_cnu_50_in_0, msg_to_check_it_2_cnu_50_in_1, msg_to_check_it_2_cnu_50_in_2, msg_to_check_it_2_cnu_50_in_3, msg_to_check_it_2_cnu_50_in_4, msg_to_check_it_2_cnu_50_in_5, msg_to_check_it_2_cnu_51_in_0, msg_to_check_it_2_cnu_51_in_1, msg_to_check_it_2_cnu_51_in_2, msg_to_check_it_2_cnu_51_in_3, msg_to_check_it_2_cnu_51_in_4, msg_to_check_it_2_cnu_51_in_5, msg_to_check_it_2_cnu_52_in_0, msg_to_check_it_2_cnu_52_in_1, msg_to_check_it_2_cnu_52_in_2, msg_to_check_it_2_cnu_52_in_3, msg_to_check_it_2_cnu_52_in_4, msg_to_check_it_2_cnu_52_in_5, msg_to_check_it_2_cnu_53_in_0, msg_to_check_it_2_cnu_53_in_1, msg_to_check_it_2_cnu_53_in_2, msg_to_check_it_2_cnu_53_in_3, msg_to_check_it_2_cnu_53_in_4, msg_to_check_it_2_cnu_53_in_5, msg_to_check_it_2_cnu_54_in_0, msg_to_check_it_2_cnu_54_in_1, msg_to_check_it_2_cnu_54_in_2, msg_to_check_it_2_cnu_54_in_3, msg_to_check_it_2_cnu_54_in_4, msg_to_check_it_2_cnu_54_in_5, msg_to_check_it_2_cnu_55_in_0, msg_to_check_it_2_cnu_55_in_1, msg_to_check_it_2_cnu_55_in_2, msg_to_check_it_2_cnu_55_in_3, msg_to_check_it_2_cnu_55_in_4, msg_to_check_it_2_cnu_55_in_5, msg_to_check_it_2_cnu_56_in_0, msg_to_check_it_2_cnu_56_in_1, msg_to_check_it_2_cnu_56_in_2, msg_to_check_it_2_cnu_56_in_3, msg_to_check_it_2_cnu_56_in_4, msg_to_check_it_2_cnu_56_in_5, msg_to_check_it_2_cnu_57_in_0, msg_to_check_it_2_cnu_57_in_1, msg_to_check_it_2_cnu_57_in_2, msg_to_check_it_2_cnu_57_in_3, msg_to_check_it_2_cnu_57_in_4, msg_to_check_it_2_cnu_57_in_5, msg_to_check_it_2_cnu_58_in_0, msg_to_check_it_2_cnu_58_in_1, msg_to_check_it_2_cnu_58_in_2, msg_to_check_it_2_cnu_58_in_3, msg_to_check_it_2_cnu_58_in_4, msg_to_check_it_2_cnu_58_in_5, msg_to_check_it_2_cnu_59_in_0, msg_to_check_it_2_cnu_59_in_1, msg_to_check_it_2_cnu_59_in_2, msg_to_check_it_2_cnu_59_in_3, msg_to_check_it_2_cnu_59_in_4, msg_to_check_it_2_cnu_59_in_5, msg_to_check_it_2_cnu_60_in_0, msg_to_check_it_2_cnu_60_in_1, msg_to_check_it_2_cnu_60_in_2, msg_to_check_it_2_cnu_60_in_3, msg_to_check_it_2_cnu_60_in_4, msg_to_check_it_2_cnu_60_in_5, msg_to_check_it_2_cnu_61_in_0, msg_to_check_it_2_cnu_61_in_1, msg_to_check_it_2_cnu_61_in_2, msg_to_check_it_2_cnu_61_in_3, msg_to_check_it_2_cnu_61_in_4, msg_to_check_it_2_cnu_61_in_5, msg_to_check_it_2_cnu_62_in_0, msg_to_check_it_2_cnu_62_in_1, msg_to_check_it_2_cnu_62_in_2, msg_to_check_it_2_cnu_62_in_3, msg_to_check_it_2_cnu_62_in_4, msg_to_check_it_2_cnu_62_in_5, msg_to_check_it_2_cnu_63_in_0, msg_to_check_it_2_cnu_63_in_1, msg_to_check_it_2_cnu_63_in_2, msg_to_check_it_2_cnu_63_in_3, msg_to_check_it_2_cnu_63_in_4, msg_to_check_it_2_cnu_63_in_5, msg_to_check_it_2_cnu_64_in_0, msg_to_check_it_2_cnu_64_in_1, msg_to_check_it_2_cnu_64_in_2, msg_to_check_it_2_cnu_64_in_3, msg_to_check_it_2_cnu_64_in_4, msg_to_check_it_2_cnu_64_in_5, msg_to_check_it_2_cnu_65_in_0, msg_to_check_it_2_cnu_65_in_1, msg_to_check_it_2_cnu_65_in_2, msg_to_check_it_2_cnu_65_in_3, msg_to_check_it_2_cnu_65_in_4, msg_to_check_it_2_cnu_65_in_5, msg_to_check_it_2_cnu_66_in_0, msg_to_check_it_2_cnu_66_in_1, msg_to_check_it_2_cnu_66_in_2, msg_to_check_it_2_cnu_66_in_3, msg_to_check_it_2_cnu_66_in_4, msg_to_check_it_2_cnu_66_in_5, msg_to_check_it_2_cnu_67_in_0, msg_to_check_it_2_cnu_67_in_1, msg_to_check_it_2_cnu_67_in_2, msg_to_check_it_2_cnu_67_in_3, msg_to_check_it_2_cnu_67_in_4, msg_to_check_it_2_cnu_67_in_5, msg_to_check_it_2_cnu_68_in_0, msg_to_check_it_2_cnu_68_in_1, msg_to_check_it_2_cnu_68_in_2, msg_to_check_it_2_cnu_68_in_3, msg_to_check_it_2_cnu_68_in_4, msg_to_check_it_2_cnu_68_in_5, msg_to_check_it_2_cnu_69_in_0, msg_to_check_it_2_cnu_69_in_1, msg_to_check_it_2_cnu_69_in_2, msg_to_check_it_2_cnu_69_in_3, msg_to_check_it_2_cnu_69_in_4, msg_to_check_it_2_cnu_69_in_5, msg_to_check_it_2_cnu_70_in_0, msg_to_check_it_2_cnu_70_in_1, msg_to_check_it_2_cnu_70_in_2, msg_to_check_it_2_cnu_70_in_3, msg_to_check_it_2_cnu_70_in_4, msg_to_check_it_2_cnu_70_in_5, msg_to_check_it_2_cnu_71_in_0, msg_to_check_it_2_cnu_71_in_1, msg_to_check_it_2_cnu_71_in_2, msg_to_check_it_2_cnu_71_in_3, msg_to_check_it_2_cnu_71_in_4, msg_to_check_it_2_cnu_71_in_5, msg_to_check_it_2_cnu_72_in_0, msg_to_check_it_2_cnu_72_in_1, msg_to_check_it_2_cnu_72_in_2, msg_to_check_it_2_cnu_72_in_3, msg_to_check_it_2_cnu_72_in_4, msg_to_check_it_2_cnu_72_in_5, msg_to_check_it_2_cnu_73_in_0, msg_to_check_it_2_cnu_73_in_1, msg_to_check_it_2_cnu_73_in_2, msg_to_check_it_2_cnu_73_in_3, msg_to_check_it_2_cnu_73_in_4, msg_to_check_it_2_cnu_73_in_5, msg_to_check_it_2_cnu_74_in_0, msg_to_check_it_2_cnu_74_in_1, msg_to_check_it_2_cnu_74_in_2, msg_to_check_it_2_cnu_74_in_3, msg_to_check_it_2_cnu_74_in_4, msg_to_check_it_2_cnu_74_in_5, msg_to_check_it_2_cnu_75_in_0, msg_to_check_it_2_cnu_75_in_1, msg_to_check_it_2_cnu_75_in_2, msg_to_check_it_2_cnu_75_in_3, msg_to_check_it_2_cnu_75_in_4, msg_to_check_it_2_cnu_75_in_5, msg_to_check_it_2_cnu_76_in_0, msg_to_check_it_2_cnu_76_in_1, msg_to_check_it_2_cnu_76_in_2, msg_to_check_it_2_cnu_76_in_3, msg_to_check_it_2_cnu_76_in_4, msg_to_check_it_2_cnu_76_in_5, msg_to_check_it_2_cnu_77_in_0, msg_to_check_it_2_cnu_77_in_1, msg_to_check_it_2_cnu_77_in_2, msg_to_check_it_2_cnu_77_in_3, msg_to_check_it_2_cnu_77_in_4, msg_to_check_it_2_cnu_77_in_5, msg_to_check_it_2_cnu_78_in_0, msg_to_check_it_2_cnu_78_in_1, msg_to_check_it_2_cnu_78_in_2, msg_to_check_it_2_cnu_78_in_3, msg_to_check_it_2_cnu_78_in_4, msg_to_check_it_2_cnu_78_in_5, msg_to_check_it_2_cnu_79_in_0, msg_to_check_it_2_cnu_79_in_1, msg_to_check_it_2_cnu_79_in_2, msg_to_check_it_2_cnu_79_in_3, msg_to_check_it_2_cnu_79_in_4, msg_to_check_it_2_cnu_79_in_5, msg_to_check_it_2_cnu_80_in_0, msg_to_check_it_2_cnu_80_in_1, msg_to_check_it_2_cnu_80_in_2, msg_to_check_it_2_cnu_80_in_3, msg_to_check_it_2_cnu_80_in_4, msg_to_check_it_2_cnu_80_in_5, msg_to_check_it_2_cnu_81_in_0, msg_to_check_it_2_cnu_81_in_1, msg_to_check_it_2_cnu_81_in_2, msg_to_check_it_2_cnu_81_in_3, msg_to_check_it_2_cnu_81_in_4, msg_to_check_it_2_cnu_81_in_5, msg_to_check_it_2_cnu_82_in_0, msg_to_check_it_2_cnu_82_in_1, msg_to_check_it_2_cnu_82_in_2, msg_to_check_it_2_cnu_82_in_3, msg_to_check_it_2_cnu_82_in_4, msg_to_check_it_2_cnu_82_in_5, msg_to_check_it_2_cnu_83_in_0, msg_to_check_it_2_cnu_83_in_1, msg_to_check_it_2_cnu_83_in_2, msg_to_check_it_2_cnu_83_in_3, msg_to_check_it_2_cnu_83_in_4, msg_to_check_it_2_cnu_83_in_5, msg_to_check_it_2_cnu_84_in_0, msg_to_check_it_2_cnu_84_in_1, msg_to_check_it_2_cnu_84_in_2, msg_to_check_it_2_cnu_84_in_3, msg_to_check_it_2_cnu_84_in_4, msg_to_check_it_2_cnu_84_in_5, msg_to_check_it_2_cnu_85_in_0, msg_to_check_it_2_cnu_85_in_1, msg_to_check_it_2_cnu_85_in_2, msg_to_check_it_2_cnu_85_in_3, msg_to_check_it_2_cnu_85_in_4, msg_to_check_it_2_cnu_85_in_5, msg_to_check_it_2_cnu_86_in_0, msg_to_check_it_2_cnu_86_in_1, msg_to_check_it_2_cnu_86_in_2, msg_to_check_it_2_cnu_86_in_3, msg_to_check_it_2_cnu_86_in_4, msg_to_check_it_2_cnu_86_in_5, msg_to_check_it_2_cnu_87_in_0, msg_to_check_it_2_cnu_87_in_1, msg_to_check_it_2_cnu_87_in_2, msg_to_check_it_2_cnu_87_in_3, msg_to_check_it_2_cnu_87_in_4, msg_to_check_it_2_cnu_87_in_5, msg_to_check_it_2_cnu_88_in_0, msg_to_check_it_2_cnu_88_in_1, msg_to_check_it_2_cnu_88_in_2, msg_to_check_it_2_cnu_88_in_3, msg_to_check_it_2_cnu_88_in_4, msg_to_check_it_2_cnu_88_in_5, msg_to_check_it_2_cnu_89_in_0, msg_to_check_it_2_cnu_89_in_1, msg_to_check_it_2_cnu_89_in_2, msg_to_check_it_2_cnu_89_in_3, msg_to_check_it_2_cnu_89_in_4, msg_to_check_it_2_cnu_89_in_5, msg_to_check_it_2_cnu_90_in_0, msg_to_check_it_2_cnu_90_in_1, msg_to_check_it_2_cnu_90_in_2, msg_to_check_it_2_cnu_90_in_3, msg_to_check_it_2_cnu_90_in_4, msg_to_check_it_2_cnu_90_in_5, msg_to_check_it_2_cnu_91_in_0, msg_to_check_it_2_cnu_91_in_1, msg_to_check_it_2_cnu_91_in_2, msg_to_check_it_2_cnu_91_in_3, msg_to_check_it_2_cnu_91_in_4, msg_to_check_it_2_cnu_91_in_5, msg_to_check_it_2_cnu_92_in_0, msg_to_check_it_2_cnu_92_in_1, msg_to_check_it_2_cnu_92_in_2, msg_to_check_it_2_cnu_92_in_3, msg_to_check_it_2_cnu_92_in_4, msg_to_check_it_2_cnu_92_in_5, msg_to_check_it_2_cnu_93_in_0, msg_to_check_it_2_cnu_93_in_1, msg_to_check_it_2_cnu_93_in_2, msg_to_check_it_2_cnu_93_in_3, msg_to_check_it_2_cnu_93_in_4, msg_to_check_it_2_cnu_93_in_5, msg_to_check_it_2_cnu_94_in_0, msg_to_check_it_2_cnu_94_in_1, msg_to_check_it_2_cnu_94_in_2, msg_to_check_it_2_cnu_94_in_3, msg_to_check_it_2_cnu_94_in_4, msg_to_check_it_2_cnu_94_in_5, msg_to_check_it_2_cnu_95_in_0, msg_to_check_it_2_cnu_95_in_1, msg_to_check_it_2_cnu_95_in_2, msg_to_check_it_2_cnu_95_in_3, msg_to_check_it_2_cnu_95_in_4, msg_to_check_it_2_cnu_95_in_5, msg_to_check_it_2_cnu_96_in_0, msg_to_check_it_2_cnu_96_in_1, msg_to_check_it_2_cnu_96_in_2, msg_to_check_it_2_cnu_96_in_3, msg_to_check_it_2_cnu_96_in_4, msg_to_check_it_2_cnu_96_in_5, msg_to_check_it_2_cnu_97_in_0, msg_to_check_it_2_cnu_97_in_1, msg_to_check_it_2_cnu_97_in_2, msg_to_check_it_2_cnu_97_in_3, msg_to_check_it_2_cnu_97_in_4, msg_to_check_it_2_cnu_97_in_5, msg_to_check_it_2_cnu_98_in_0, msg_to_check_it_2_cnu_98_in_1, msg_to_check_it_2_cnu_98_in_2, msg_to_check_it_2_cnu_98_in_3, msg_to_check_it_2_cnu_98_in_4, msg_to_check_it_2_cnu_98_in_5, msg_to_check_it_3_cnu_0_in_0, msg_to_check_it_3_cnu_0_in_1, msg_to_check_it_3_cnu_0_in_2, msg_to_check_it_3_cnu_0_in_3, msg_to_check_it_3_cnu_0_in_4, msg_to_check_it_3_cnu_0_in_5, msg_to_check_it_3_cnu_1_in_0, msg_to_check_it_3_cnu_1_in_1, msg_to_check_it_3_cnu_1_in_2, msg_to_check_it_3_cnu_1_in_3, msg_to_check_it_3_cnu_1_in_4, msg_to_check_it_3_cnu_1_in_5, msg_to_check_it_3_cnu_2_in_0, msg_to_check_it_3_cnu_2_in_1, msg_to_check_it_3_cnu_2_in_2, msg_to_check_it_3_cnu_2_in_3, msg_to_check_it_3_cnu_2_in_4, msg_to_check_it_3_cnu_2_in_5, msg_to_check_it_3_cnu_3_in_0, msg_to_check_it_3_cnu_3_in_1, msg_to_check_it_3_cnu_3_in_2, msg_to_check_it_3_cnu_3_in_3, msg_to_check_it_3_cnu_3_in_4, msg_to_check_it_3_cnu_3_in_5, msg_to_check_it_3_cnu_4_in_0, msg_to_check_it_3_cnu_4_in_1, msg_to_check_it_3_cnu_4_in_2, msg_to_check_it_3_cnu_4_in_3, msg_to_check_it_3_cnu_4_in_4, msg_to_check_it_3_cnu_4_in_5, msg_to_check_it_3_cnu_5_in_0, msg_to_check_it_3_cnu_5_in_1, msg_to_check_it_3_cnu_5_in_2, msg_to_check_it_3_cnu_5_in_3, msg_to_check_it_3_cnu_5_in_4, msg_to_check_it_3_cnu_5_in_5, msg_to_check_it_3_cnu_6_in_0, msg_to_check_it_3_cnu_6_in_1, msg_to_check_it_3_cnu_6_in_2, msg_to_check_it_3_cnu_6_in_3, msg_to_check_it_3_cnu_6_in_4, msg_to_check_it_3_cnu_6_in_5, msg_to_check_it_3_cnu_7_in_0, msg_to_check_it_3_cnu_7_in_1, msg_to_check_it_3_cnu_7_in_2, msg_to_check_it_3_cnu_7_in_3, msg_to_check_it_3_cnu_7_in_4, msg_to_check_it_3_cnu_7_in_5, msg_to_check_it_3_cnu_8_in_0, msg_to_check_it_3_cnu_8_in_1, msg_to_check_it_3_cnu_8_in_2, msg_to_check_it_3_cnu_8_in_3, msg_to_check_it_3_cnu_8_in_4, msg_to_check_it_3_cnu_8_in_5, msg_to_check_it_3_cnu_9_in_0, msg_to_check_it_3_cnu_9_in_1, msg_to_check_it_3_cnu_9_in_2, msg_to_check_it_3_cnu_9_in_3, msg_to_check_it_3_cnu_9_in_4, msg_to_check_it_3_cnu_9_in_5, msg_to_check_it_3_cnu_10_in_0, msg_to_check_it_3_cnu_10_in_1, msg_to_check_it_3_cnu_10_in_2, msg_to_check_it_3_cnu_10_in_3, msg_to_check_it_3_cnu_10_in_4, msg_to_check_it_3_cnu_10_in_5, msg_to_check_it_3_cnu_11_in_0, msg_to_check_it_3_cnu_11_in_1, msg_to_check_it_3_cnu_11_in_2, msg_to_check_it_3_cnu_11_in_3, msg_to_check_it_3_cnu_11_in_4, msg_to_check_it_3_cnu_11_in_5, msg_to_check_it_3_cnu_12_in_0, msg_to_check_it_3_cnu_12_in_1, msg_to_check_it_3_cnu_12_in_2, msg_to_check_it_3_cnu_12_in_3, msg_to_check_it_3_cnu_12_in_4, msg_to_check_it_3_cnu_12_in_5, msg_to_check_it_3_cnu_13_in_0, msg_to_check_it_3_cnu_13_in_1, msg_to_check_it_3_cnu_13_in_2, msg_to_check_it_3_cnu_13_in_3, msg_to_check_it_3_cnu_13_in_4, msg_to_check_it_3_cnu_13_in_5, msg_to_check_it_3_cnu_14_in_0, msg_to_check_it_3_cnu_14_in_1, msg_to_check_it_3_cnu_14_in_2, msg_to_check_it_3_cnu_14_in_3, msg_to_check_it_3_cnu_14_in_4, msg_to_check_it_3_cnu_14_in_5, msg_to_check_it_3_cnu_15_in_0, msg_to_check_it_3_cnu_15_in_1, msg_to_check_it_3_cnu_15_in_2, msg_to_check_it_3_cnu_15_in_3, msg_to_check_it_3_cnu_15_in_4, msg_to_check_it_3_cnu_15_in_5, msg_to_check_it_3_cnu_16_in_0, msg_to_check_it_3_cnu_16_in_1, msg_to_check_it_3_cnu_16_in_2, msg_to_check_it_3_cnu_16_in_3, msg_to_check_it_3_cnu_16_in_4, msg_to_check_it_3_cnu_16_in_5, msg_to_check_it_3_cnu_17_in_0, msg_to_check_it_3_cnu_17_in_1, msg_to_check_it_3_cnu_17_in_2, msg_to_check_it_3_cnu_17_in_3, msg_to_check_it_3_cnu_17_in_4, msg_to_check_it_3_cnu_17_in_5, msg_to_check_it_3_cnu_18_in_0, msg_to_check_it_3_cnu_18_in_1, msg_to_check_it_3_cnu_18_in_2, msg_to_check_it_3_cnu_18_in_3, msg_to_check_it_3_cnu_18_in_4, msg_to_check_it_3_cnu_18_in_5, msg_to_check_it_3_cnu_19_in_0, msg_to_check_it_3_cnu_19_in_1, msg_to_check_it_3_cnu_19_in_2, msg_to_check_it_3_cnu_19_in_3, msg_to_check_it_3_cnu_19_in_4, msg_to_check_it_3_cnu_19_in_5, msg_to_check_it_3_cnu_20_in_0, msg_to_check_it_3_cnu_20_in_1, msg_to_check_it_3_cnu_20_in_2, msg_to_check_it_3_cnu_20_in_3, msg_to_check_it_3_cnu_20_in_4, msg_to_check_it_3_cnu_20_in_5, msg_to_check_it_3_cnu_21_in_0, msg_to_check_it_3_cnu_21_in_1, msg_to_check_it_3_cnu_21_in_2, msg_to_check_it_3_cnu_21_in_3, msg_to_check_it_3_cnu_21_in_4, msg_to_check_it_3_cnu_21_in_5, msg_to_check_it_3_cnu_22_in_0, msg_to_check_it_3_cnu_22_in_1, msg_to_check_it_3_cnu_22_in_2, msg_to_check_it_3_cnu_22_in_3, msg_to_check_it_3_cnu_22_in_4, msg_to_check_it_3_cnu_22_in_5, msg_to_check_it_3_cnu_23_in_0, msg_to_check_it_3_cnu_23_in_1, msg_to_check_it_3_cnu_23_in_2, msg_to_check_it_3_cnu_23_in_3, msg_to_check_it_3_cnu_23_in_4, msg_to_check_it_3_cnu_23_in_5, msg_to_check_it_3_cnu_24_in_0, msg_to_check_it_3_cnu_24_in_1, msg_to_check_it_3_cnu_24_in_2, msg_to_check_it_3_cnu_24_in_3, msg_to_check_it_3_cnu_24_in_4, msg_to_check_it_3_cnu_24_in_5, msg_to_check_it_3_cnu_25_in_0, msg_to_check_it_3_cnu_25_in_1, msg_to_check_it_3_cnu_25_in_2, msg_to_check_it_3_cnu_25_in_3, msg_to_check_it_3_cnu_25_in_4, msg_to_check_it_3_cnu_25_in_5, msg_to_check_it_3_cnu_26_in_0, msg_to_check_it_3_cnu_26_in_1, msg_to_check_it_3_cnu_26_in_2, msg_to_check_it_3_cnu_26_in_3, msg_to_check_it_3_cnu_26_in_4, msg_to_check_it_3_cnu_26_in_5, msg_to_check_it_3_cnu_27_in_0, msg_to_check_it_3_cnu_27_in_1, msg_to_check_it_3_cnu_27_in_2, msg_to_check_it_3_cnu_27_in_3, msg_to_check_it_3_cnu_27_in_4, msg_to_check_it_3_cnu_27_in_5, msg_to_check_it_3_cnu_28_in_0, msg_to_check_it_3_cnu_28_in_1, msg_to_check_it_3_cnu_28_in_2, msg_to_check_it_3_cnu_28_in_3, msg_to_check_it_3_cnu_28_in_4, msg_to_check_it_3_cnu_28_in_5, msg_to_check_it_3_cnu_29_in_0, msg_to_check_it_3_cnu_29_in_1, msg_to_check_it_3_cnu_29_in_2, msg_to_check_it_3_cnu_29_in_3, msg_to_check_it_3_cnu_29_in_4, msg_to_check_it_3_cnu_29_in_5, msg_to_check_it_3_cnu_30_in_0, msg_to_check_it_3_cnu_30_in_1, msg_to_check_it_3_cnu_30_in_2, msg_to_check_it_3_cnu_30_in_3, msg_to_check_it_3_cnu_30_in_4, msg_to_check_it_3_cnu_30_in_5, msg_to_check_it_3_cnu_31_in_0, msg_to_check_it_3_cnu_31_in_1, msg_to_check_it_3_cnu_31_in_2, msg_to_check_it_3_cnu_31_in_3, msg_to_check_it_3_cnu_31_in_4, msg_to_check_it_3_cnu_31_in_5, msg_to_check_it_3_cnu_32_in_0, msg_to_check_it_3_cnu_32_in_1, msg_to_check_it_3_cnu_32_in_2, msg_to_check_it_3_cnu_32_in_3, msg_to_check_it_3_cnu_32_in_4, msg_to_check_it_3_cnu_32_in_5, msg_to_check_it_3_cnu_33_in_0, msg_to_check_it_3_cnu_33_in_1, msg_to_check_it_3_cnu_33_in_2, msg_to_check_it_3_cnu_33_in_3, msg_to_check_it_3_cnu_33_in_4, msg_to_check_it_3_cnu_33_in_5, msg_to_check_it_3_cnu_34_in_0, msg_to_check_it_3_cnu_34_in_1, msg_to_check_it_3_cnu_34_in_2, msg_to_check_it_3_cnu_34_in_3, msg_to_check_it_3_cnu_34_in_4, msg_to_check_it_3_cnu_34_in_5, msg_to_check_it_3_cnu_35_in_0, msg_to_check_it_3_cnu_35_in_1, msg_to_check_it_3_cnu_35_in_2, msg_to_check_it_3_cnu_35_in_3, msg_to_check_it_3_cnu_35_in_4, msg_to_check_it_3_cnu_35_in_5, msg_to_check_it_3_cnu_36_in_0, msg_to_check_it_3_cnu_36_in_1, msg_to_check_it_3_cnu_36_in_2, msg_to_check_it_3_cnu_36_in_3, msg_to_check_it_3_cnu_36_in_4, msg_to_check_it_3_cnu_36_in_5, msg_to_check_it_3_cnu_37_in_0, msg_to_check_it_3_cnu_37_in_1, msg_to_check_it_3_cnu_37_in_2, msg_to_check_it_3_cnu_37_in_3, msg_to_check_it_3_cnu_37_in_4, msg_to_check_it_3_cnu_37_in_5, msg_to_check_it_3_cnu_38_in_0, msg_to_check_it_3_cnu_38_in_1, msg_to_check_it_3_cnu_38_in_2, msg_to_check_it_3_cnu_38_in_3, msg_to_check_it_3_cnu_38_in_4, msg_to_check_it_3_cnu_38_in_5, msg_to_check_it_3_cnu_39_in_0, msg_to_check_it_3_cnu_39_in_1, msg_to_check_it_3_cnu_39_in_2, msg_to_check_it_3_cnu_39_in_3, msg_to_check_it_3_cnu_39_in_4, msg_to_check_it_3_cnu_39_in_5, msg_to_check_it_3_cnu_40_in_0, msg_to_check_it_3_cnu_40_in_1, msg_to_check_it_3_cnu_40_in_2, msg_to_check_it_3_cnu_40_in_3, msg_to_check_it_3_cnu_40_in_4, msg_to_check_it_3_cnu_40_in_5, msg_to_check_it_3_cnu_41_in_0, msg_to_check_it_3_cnu_41_in_1, msg_to_check_it_3_cnu_41_in_2, msg_to_check_it_3_cnu_41_in_3, msg_to_check_it_3_cnu_41_in_4, msg_to_check_it_3_cnu_41_in_5, msg_to_check_it_3_cnu_42_in_0, msg_to_check_it_3_cnu_42_in_1, msg_to_check_it_3_cnu_42_in_2, msg_to_check_it_3_cnu_42_in_3, msg_to_check_it_3_cnu_42_in_4, msg_to_check_it_3_cnu_42_in_5, msg_to_check_it_3_cnu_43_in_0, msg_to_check_it_3_cnu_43_in_1, msg_to_check_it_3_cnu_43_in_2, msg_to_check_it_3_cnu_43_in_3, msg_to_check_it_3_cnu_43_in_4, msg_to_check_it_3_cnu_43_in_5, msg_to_check_it_3_cnu_44_in_0, msg_to_check_it_3_cnu_44_in_1, msg_to_check_it_3_cnu_44_in_2, msg_to_check_it_3_cnu_44_in_3, msg_to_check_it_3_cnu_44_in_4, msg_to_check_it_3_cnu_44_in_5, msg_to_check_it_3_cnu_45_in_0, msg_to_check_it_3_cnu_45_in_1, msg_to_check_it_3_cnu_45_in_2, msg_to_check_it_3_cnu_45_in_3, msg_to_check_it_3_cnu_45_in_4, msg_to_check_it_3_cnu_45_in_5, msg_to_check_it_3_cnu_46_in_0, msg_to_check_it_3_cnu_46_in_1, msg_to_check_it_3_cnu_46_in_2, msg_to_check_it_3_cnu_46_in_3, msg_to_check_it_3_cnu_46_in_4, msg_to_check_it_3_cnu_46_in_5, msg_to_check_it_3_cnu_47_in_0, msg_to_check_it_3_cnu_47_in_1, msg_to_check_it_3_cnu_47_in_2, msg_to_check_it_3_cnu_47_in_3, msg_to_check_it_3_cnu_47_in_4, msg_to_check_it_3_cnu_47_in_5, msg_to_check_it_3_cnu_48_in_0, msg_to_check_it_3_cnu_48_in_1, msg_to_check_it_3_cnu_48_in_2, msg_to_check_it_3_cnu_48_in_3, msg_to_check_it_3_cnu_48_in_4, msg_to_check_it_3_cnu_48_in_5, msg_to_check_it_3_cnu_49_in_0, msg_to_check_it_3_cnu_49_in_1, msg_to_check_it_3_cnu_49_in_2, msg_to_check_it_3_cnu_49_in_3, msg_to_check_it_3_cnu_49_in_4, msg_to_check_it_3_cnu_49_in_5, msg_to_check_it_3_cnu_50_in_0, msg_to_check_it_3_cnu_50_in_1, msg_to_check_it_3_cnu_50_in_2, msg_to_check_it_3_cnu_50_in_3, msg_to_check_it_3_cnu_50_in_4, msg_to_check_it_3_cnu_50_in_5, msg_to_check_it_3_cnu_51_in_0, msg_to_check_it_3_cnu_51_in_1, msg_to_check_it_3_cnu_51_in_2, msg_to_check_it_3_cnu_51_in_3, msg_to_check_it_3_cnu_51_in_4, msg_to_check_it_3_cnu_51_in_5, msg_to_check_it_3_cnu_52_in_0, msg_to_check_it_3_cnu_52_in_1, msg_to_check_it_3_cnu_52_in_2, msg_to_check_it_3_cnu_52_in_3, msg_to_check_it_3_cnu_52_in_4, msg_to_check_it_3_cnu_52_in_5, msg_to_check_it_3_cnu_53_in_0, msg_to_check_it_3_cnu_53_in_1, msg_to_check_it_3_cnu_53_in_2, msg_to_check_it_3_cnu_53_in_3, msg_to_check_it_3_cnu_53_in_4, msg_to_check_it_3_cnu_53_in_5, msg_to_check_it_3_cnu_54_in_0, msg_to_check_it_3_cnu_54_in_1, msg_to_check_it_3_cnu_54_in_2, msg_to_check_it_3_cnu_54_in_3, msg_to_check_it_3_cnu_54_in_4, msg_to_check_it_3_cnu_54_in_5, msg_to_check_it_3_cnu_55_in_0, msg_to_check_it_3_cnu_55_in_1, msg_to_check_it_3_cnu_55_in_2, msg_to_check_it_3_cnu_55_in_3, msg_to_check_it_3_cnu_55_in_4, msg_to_check_it_3_cnu_55_in_5, msg_to_check_it_3_cnu_56_in_0, msg_to_check_it_3_cnu_56_in_1, msg_to_check_it_3_cnu_56_in_2, msg_to_check_it_3_cnu_56_in_3, msg_to_check_it_3_cnu_56_in_4, msg_to_check_it_3_cnu_56_in_5, msg_to_check_it_3_cnu_57_in_0, msg_to_check_it_3_cnu_57_in_1, msg_to_check_it_3_cnu_57_in_2, msg_to_check_it_3_cnu_57_in_3, msg_to_check_it_3_cnu_57_in_4, msg_to_check_it_3_cnu_57_in_5, msg_to_check_it_3_cnu_58_in_0, msg_to_check_it_3_cnu_58_in_1, msg_to_check_it_3_cnu_58_in_2, msg_to_check_it_3_cnu_58_in_3, msg_to_check_it_3_cnu_58_in_4, msg_to_check_it_3_cnu_58_in_5, msg_to_check_it_3_cnu_59_in_0, msg_to_check_it_3_cnu_59_in_1, msg_to_check_it_3_cnu_59_in_2, msg_to_check_it_3_cnu_59_in_3, msg_to_check_it_3_cnu_59_in_4, msg_to_check_it_3_cnu_59_in_5, msg_to_check_it_3_cnu_60_in_0, msg_to_check_it_3_cnu_60_in_1, msg_to_check_it_3_cnu_60_in_2, msg_to_check_it_3_cnu_60_in_3, msg_to_check_it_3_cnu_60_in_4, msg_to_check_it_3_cnu_60_in_5, msg_to_check_it_3_cnu_61_in_0, msg_to_check_it_3_cnu_61_in_1, msg_to_check_it_3_cnu_61_in_2, msg_to_check_it_3_cnu_61_in_3, msg_to_check_it_3_cnu_61_in_4, msg_to_check_it_3_cnu_61_in_5, msg_to_check_it_3_cnu_62_in_0, msg_to_check_it_3_cnu_62_in_1, msg_to_check_it_3_cnu_62_in_2, msg_to_check_it_3_cnu_62_in_3, msg_to_check_it_3_cnu_62_in_4, msg_to_check_it_3_cnu_62_in_5, msg_to_check_it_3_cnu_63_in_0, msg_to_check_it_3_cnu_63_in_1, msg_to_check_it_3_cnu_63_in_2, msg_to_check_it_3_cnu_63_in_3, msg_to_check_it_3_cnu_63_in_4, msg_to_check_it_3_cnu_63_in_5, msg_to_check_it_3_cnu_64_in_0, msg_to_check_it_3_cnu_64_in_1, msg_to_check_it_3_cnu_64_in_2, msg_to_check_it_3_cnu_64_in_3, msg_to_check_it_3_cnu_64_in_4, msg_to_check_it_3_cnu_64_in_5, msg_to_check_it_3_cnu_65_in_0, msg_to_check_it_3_cnu_65_in_1, msg_to_check_it_3_cnu_65_in_2, msg_to_check_it_3_cnu_65_in_3, msg_to_check_it_3_cnu_65_in_4, msg_to_check_it_3_cnu_65_in_5, msg_to_check_it_3_cnu_66_in_0, msg_to_check_it_3_cnu_66_in_1, msg_to_check_it_3_cnu_66_in_2, msg_to_check_it_3_cnu_66_in_3, msg_to_check_it_3_cnu_66_in_4, msg_to_check_it_3_cnu_66_in_5, msg_to_check_it_3_cnu_67_in_0, msg_to_check_it_3_cnu_67_in_1, msg_to_check_it_3_cnu_67_in_2, msg_to_check_it_3_cnu_67_in_3, msg_to_check_it_3_cnu_67_in_4, msg_to_check_it_3_cnu_67_in_5, msg_to_check_it_3_cnu_68_in_0, msg_to_check_it_3_cnu_68_in_1, msg_to_check_it_3_cnu_68_in_2, msg_to_check_it_3_cnu_68_in_3, msg_to_check_it_3_cnu_68_in_4, msg_to_check_it_3_cnu_68_in_5, msg_to_check_it_3_cnu_69_in_0, msg_to_check_it_3_cnu_69_in_1, msg_to_check_it_3_cnu_69_in_2, msg_to_check_it_3_cnu_69_in_3, msg_to_check_it_3_cnu_69_in_4, msg_to_check_it_3_cnu_69_in_5, msg_to_check_it_3_cnu_70_in_0, msg_to_check_it_3_cnu_70_in_1, msg_to_check_it_3_cnu_70_in_2, msg_to_check_it_3_cnu_70_in_3, msg_to_check_it_3_cnu_70_in_4, msg_to_check_it_3_cnu_70_in_5, msg_to_check_it_3_cnu_71_in_0, msg_to_check_it_3_cnu_71_in_1, msg_to_check_it_3_cnu_71_in_2, msg_to_check_it_3_cnu_71_in_3, msg_to_check_it_3_cnu_71_in_4, msg_to_check_it_3_cnu_71_in_5, msg_to_check_it_3_cnu_72_in_0, msg_to_check_it_3_cnu_72_in_1, msg_to_check_it_3_cnu_72_in_2, msg_to_check_it_3_cnu_72_in_3, msg_to_check_it_3_cnu_72_in_4, msg_to_check_it_3_cnu_72_in_5, msg_to_check_it_3_cnu_73_in_0, msg_to_check_it_3_cnu_73_in_1, msg_to_check_it_3_cnu_73_in_2, msg_to_check_it_3_cnu_73_in_3, msg_to_check_it_3_cnu_73_in_4, msg_to_check_it_3_cnu_73_in_5, msg_to_check_it_3_cnu_74_in_0, msg_to_check_it_3_cnu_74_in_1, msg_to_check_it_3_cnu_74_in_2, msg_to_check_it_3_cnu_74_in_3, msg_to_check_it_3_cnu_74_in_4, msg_to_check_it_3_cnu_74_in_5, msg_to_check_it_3_cnu_75_in_0, msg_to_check_it_3_cnu_75_in_1, msg_to_check_it_3_cnu_75_in_2, msg_to_check_it_3_cnu_75_in_3, msg_to_check_it_3_cnu_75_in_4, msg_to_check_it_3_cnu_75_in_5, msg_to_check_it_3_cnu_76_in_0, msg_to_check_it_3_cnu_76_in_1, msg_to_check_it_3_cnu_76_in_2, msg_to_check_it_3_cnu_76_in_3, msg_to_check_it_3_cnu_76_in_4, msg_to_check_it_3_cnu_76_in_5, msg_to_check_it_3_cnu_77_in_0, msg_to_check_it_3_cnu_77_in_1, msg_to_check_it_3_cnu_77_in_2, msg_to_check_it_3_cnu_77_in_3, msg_to_check_it_3_cnu_77_in_4, msg_to_check_it_3_cnu_77_in_5, msg_to_check_it_3_cnu_78_in_0, msg_to_check_it_3_cnu_78_in_1, msg_to_check_it_3_cnu_78_in_2, msg_to_check_it_3_cnu_78_in_3, msg_to_check_it_3_cnu_78_in_4, msg_to_check_it_3_cnu_78_in_5, msg_to_check_it_3_cnu_79_in_0, msg_to_check_it_3_cnu_79_in_1, msg_to_check_it_3_cnu_79_in_2, msg_to_check_it_3_cnu_79_in_3, msg_to_check_it_3_cnu_79_in_4, msg_to_check_it_3_cnu_79_in_5, msg_to_check_it_3_cnu_80_in_0, msg_to_check_it_3_cnu_80_in_1, msg_to_check_it_3_cnu_80_in_2, msg_to_check_it_3_cnu_80_in_3, msg_to_check_it_3_cnu_80_in_4, msg_to_check_it_3_cnu_80_in_5, msg_to_check_it_3_cnu_81_in_0, msg_to_check_it_3_cnu_81_in_1, msg_to_check_it_3_cnu_81_in_2, msg_to_check_it_3_cnu_81_in_3, msg_to_check_it_3_cnu_81_in_4, msg_to_check_it_3_cnu_81_in_5, msg_to_check_it_3_cnu_82_in_0, msg_to_check_it_3_cnu_82_in_1, msg_to_check_it_3_cnu_82_in_2, msg_to_check_it_3_cnu_82_in_3, msg_to_check_it_3_cnu_82_in_4, msg_to_check_it_3_cnu_82_in_5, msg_to_check_it_3_cnu_83_in_0, msg_to_check_it_3_cnu_83_in_1, msg_to_check_it_3_cnu_83_in_2, msg_to_check_it_3_cnu_83_in_3, msg_to_check_it_3_cnu_83_in_4, msg_to_check_it_3_cnu_83_in_5, msg_to_check_it_3_cnu_84_in_0, msg_to_check_it_3_cnu_84_in_1, msg_to_check_it_3_cnu_84_in_2, msg_to_check_it_3_cnu_84_in_3, msg_to_check_it_3_cnu_84_in_4, msg_to_check_it_3_cnu_84_in_5, msg_to_check_it_3_cnu_85_in_0, msg_to_check_it_3_cnu_85_in_1, msg_to_check_it_3_cnu_85_in_2, msg_to_check_it_3_cnu_85_in_3, msg_to_check_it_3_cnu_85_in_4, msg_to_check_it_3_cnu_85_in_5, msg_to_check_it_3_cnu_86_in_0, msg_to_check_it_3_cnu_86_in_1, msg_to_check_it_3_cnu_86_in_2, msg_to_check_it_3_cnu_86_in_3, msg_to_check_it_3_cnu_86_in_4, msg_to_check_it_3_cnu_86_in_5, msg_to_check_it_3_cnu_87_in_0, msg_to_check_it_3_cnu_87_in_1, msg_to_check_it_3_cnu_87_in_2, msg_to_check_it_3_cnu_87_in_3, msg_to_check_it_3_cnu_87_in_4, msg_to_check_it_3_cnu_87_in_5, msg_to_check_it_3_cnu_88_in_0, msg_to_check_it_3_cnu_88_in_1, msg_to_check_it_3_cnu_88_in_2, msg_to_check_it_3_cnu_88_in_3, msg_to_check_it_3_cnu_88_in_4, msg_to_check_it_3_cnu_88_in_5, msg_to_check_it_3_cnu_89_in_0, msg_to_check_it_3_cnu_89_in_1, msg_to_check_it_3_cnu_89_in_2, msg_to_check_it_3_cnu_89_in_3, msg_to_check_it_3_cnu_89_in_4, msg_to_check_it_3_cnu_89_in_5, msg_to_check_it_3_cnu_90_in_0, msg_to_check_it_3_cnu_90_in_1, msg_to_check_it_3_cnu_90_in_2, msg_to_check_it_3_cnu_90_in_3, msg_to_check_it_3_cnu_90_in_4, msg_to_check_it_3_cnu_90_in_5, msg_to_check_it_3_cnu_91_in_0, msg_to_check_it_3_cnu_91_in_1, msg_to_check_it_3_cnu_91_in_2, msg_to_check_it_3_cnu_91_in_3, msg_to_check_it_3_cnu_91_in_4, msg_to_check_it_3_cnu_91_in_5, msg_to_check_it_3_cnu_92_in_0, msg_to_check_it_3_cnu_92_in_1, msg_to_check_it_3_cnu_92_in_2, msg_to_check_it_3_cnu_92_in_3, msg_to_check_it_3_cnu_92_in_4, msg_to_check_it_3_cnu_92_in_5, msg_to_check_it_3_cnu_93_in_0, msg_to_check_it_3_cnu_93_in_1, msg_to_check_it_3_cnu_93_in_2, msg_to_check_it_3_cnu_93_in_3, msg_to_check_it_3_cnu_93_in_4, msg_to_check_it_3_cnu_93_in_5, msg_to_check_it_3_cnu_94_in_0, msg_to_check_it_3_cnu_94_in_1, msg_to_check_it_3_cnu_94_in_2, msg_to_check_it_3_cnu_94_in_3, msg_to_check_it_3_cnu_94_in_4, msg_to_check_it_3_cnu_94_in_5, msg_to_check_it_3_cnu_95_in_0, msg_to_check_it_3_cnu_95_in_1, msg_to_check_it_3_cnu_95_in_2, msg_to_check_it_3_cnu_95_in_3, msg_to_check_it_3_cnu_95_in_4, msg_to_check_it_3_cnu_95_in_5, msg_to_check_it_3_cnu_96_in_0, msg_to_check_it_3_cnu_96_in_1, msg_to_check_it_3_cnu_96_in_2, msg_to_check_it_3_cnu_96_in_3, msg_to_check_it_3_cnu_96_in_4, msg_to_check_it_3_cnu_96_in_5, msg_to_check_it_3_cnu_97_in_0, msg_to_check_it_3_cnu_97_in_1, msg_to_check_it_3_cnu_97_in_2, msg_to_check_it_3_cnu_97_in_3, msg_to_check_it_3_cnu_97_in_4, msg_to_check_it_3_cnu_97_in_5, msg_to_check_it_3_cnu_98_in_0, msg_to_check_it_3_cnu_98_in_1, msg_to_check_it_3_cnu_98_in_2, msg_to_check_it_3_cnu_98_in_3, msg_to_check_it_3_cnu_98_in_4, msg_to_check_it_3_cnu_98_in_5, msg_to_check_it_4_cnu_0_in_0, msg_to_check_it_4_cnu_0_in_1, msg_to_check_it_4_cnu_0_in_2, msg_to_check_it_4_cnu_0_in_3, msg_to_check_it_4_cnu_0_in_4, msg_to_check_it_4_cnu_0_in_5, msg_to_check_it_4_cnu_1_in_0, msg_to_check_it_4_cnu_1_in_1, msg_to_check_it_4_cnu_1_in_2, msg_to_check_it_4_cnu_1_in_3, msg_to_check_it_4_cnu_1_in_4, msg_to_check_it_4_cnu_1_in_5, msg_to_check_it_4_cnu_2_in_0, msg_to_check_it_4_cnu_2_in_1, msg_to_check_it_4_cnu_2_in_2, msg_to_check_it_4_cnu_2_in_3, msg_to_check_it_4_cnu_2_in_4, msg_to_check_it_4_cnu_2_in_5, msg_to_check_it_4_cnu_3_in_0, msg_to_check_it_4_cnu_3_in_1, msg_to_check_it_4_cnu_3_in_2, msg_to_check_it_4_cnu_3_in_3, msg_to_check_it_4_cnu_3_in_4, msg_to_check_it_4_cnu_3_in_5, msg_to_check_it_4_cnu_4_in_0, msg_to_check_it_4_cnu_4_in_1, msg_to_check_it_4_cnu_4_in_2, msg_to_check_it_4_cnu_4_in_3, msg_to_check_it_4_cnu_4_in_4, msg_to_check_it_4_cnu_4_in_5, msg_to_check_it_4_cnu_5_in_0, msg_to_check_it_4_cnu_5_in_1, msg_to_check_it_4_cnu_5_in_2, msg_to_check_it_4_cnu_5_in_3, msg_to_check_it_4_cnu_5_in_4, msg_to_check_it_4_cnu_5_in_5, msg_to_check_it_4_cnu_6_in_0, msg_to_check_it_4_cnu_6_in_1, msg_to_check_it_4_cnu_6_in_2, msg_to_check_it_4_cnu_6_in_3, msg_to_check_it_4_cnu_6_in_4, msg_to_check_it_4_cnu_6_in_5, msg_to_check_it_4_cnu_7_in_0, msg_to_check_it_4_cnu_7_in_1, msg_to_check_it_4_cnu_7_in_2, msg_to_check_it_4_cnu_7_in_3, msg_to_check_it_4_cnu_7_in_4, msg_to_check_it_4_cnu_7_in_5, msg_to_check_it_4_cnu_8_in_0, msg_to_check_it_4_cnu_8_in_1, msg_to_check_it_4_cnu_8_in_2, msg_to_check_it_4_cnu_8_in_3, msg_to_check_it_4_cnu_8_in_4, msg_to_check_it_4_cnu_8_in_5, msg_to_check_it_4_cnu_9_in_0, msg_to_check_it_4_cnu_9_in_1, msg_to_check_it_4_cnu_9_in_2, msg_to_check_it_4_cnu_9_in_3, msg_to_check_it_4_cnu_9_in_4, msg_to_check_it_4_cnu_9_in_5, msg_to_check_it_4_cnu_10_in_0, msg_to_check_it_4_cnu_10_in_1, msg_to_check_it_4_cnu_10_in_2, msg_to_check_it_4_cnu_10_in_3, msg_to_check_it_4_cnu_10_in_4, msg_to_check_it_4_cnu_10_in_5, msg_to_check_it_4_cnu_11_in_0, msg_to_check_it_4_cnu_11_in_1, msg_to_check_it_4_cnu_11_in_2, msg_to_check_it_4_cnu_11_in_3, msg_to_check_it_4_cnu_11_in_4, msg_to_check_it_4_cnu_11_in_5, msg_to_check_it_4_cnu_12_in_0, msg_to_check_it_4_cnu_12_in_1, msg_to_check_it_4_cnu_12_in_2, msg_to_check_it_4_cnu_12_in_3, msg_to_check_it_4_cnu_12_in_4, msg_to_check_it_4_cnu_12_in_5, msg_to_check_it_4_cnu_13_in_0, msg_to_check_it_4_cnu_13_in_1, msg_to_check_it_4_cnu_13_in_2, msg_to_check_it_4_cnu_13_in_3, msg_to_check_it_4_cnu_13_in_4, msg_to_check_it_4_cnu_13_in_5, msg_to_check_it_4_cnu_14_in_0, msg_to_check_it_4_cnu_14_in_1, msg_to_check_it_4_cnu_14_in_2, msg_to_check_it_4_cnu_14_in_3, msg_to_check_it_4_cnu_14_in_4, msg_to_check_it_4_cnu_14_in_5, msg_to_check_it_4_cnu_15_in_0, msg_to_check_it_4_cnu_15_in_1, msg_to_check_it_4_cnu_15_in_2, msg_to_check_it_4_cnu_15_in_3, msg_to_check_it_4_cnu_15_in_4, msg_to_check_it_4_cnu_15_in_5, msg_to_check_it_4_cnu_16_in_0, msg_to_check_it_4_cnu_16_in_1, msg_to_check_it_4_cnu_16_in_2, msg_to_check_it_4_cnu_16_in_3, msg_to_check_it_4_cnu_16_in_4, msg_to_check_it_4_cnu_16_in_5, msg_to_check_it_4_cnu_17_in_0, msg_to_check_it_4_cnu_17_in_1, msg_to_check_it_4_cnu_17_in_2, msg_to_check_it_4_cnu_17_in_3, msg_to_check_it_4_cnu_17_in_4, msg_to_check_it_4_cnu_17_in_5, msg_to_check_it_4_cnu_18_in_0, msg_to_check_it_4_cnu_18_in_1, msg_to_check_it_4_cnu_18_in_2, msg_to_check_it_4_cnu_18_in_3, msg_to_check_it_4_cnu_18_in_4, msg_to_check_it_4_cnu_18_in_5, msg_to_check_it_4_cnu_19_in_0, msg_to_check_it_4_cnu_19_in_1, msg_to_check_it_4_cnu_19_in_2, msg_to_check_it_4_cnu_19_in_3, msg_to_check_it_4_cnu_19_in_4, msg_to_check_it_4_cnu_19_in_5, msg_to_check_it_4_cnu_20_in_0, msg_to_check_it_4_cnu_20_in_1, msg_to_check_it_4_cnu_20_in_2, msg_to_check_it_4_cnu_20_in_3, msg_to_check_it_4_cnu_20_in_4, msg_to_check_it_4_cnu_20_in_5, msg_to_check_it_4_cnu_21_in_0, msg_to_check_it_4_cnu_21_in_1, msg_to_check_it_4_cnu_21_in_2, msg_to_check_it_4_cnu_21_in_3, msg_to_check_it_4_cnu_21_in_4, msg_to_check_it_4_cnu_21_in_5, msg_to_check_it_4_cnu_22_in_0, msg_to_check_it_4_cnu_22_in_1, msg_to_check_it_4_cnu_22_in_2, msg_to_check_it_4_cnu_22_in_3, msg_to_check_it_4_cnu_22_in_4, msg_to_check_it_4_cnu_22_in_5, msg_to_check_it_4_cnu_23_in_0, msg_to_check_it_4_cnu_23_in_1, msg_to_check_it_4_cnu_23_in_2, msg_to_check_it_4_cnu_23_in_3, msg_to_check_it_4_cnu_23_in_4, msg_to_check_it_4_cnu_23_in_5, msg_to_check_it_4_cnu_24_in_0, msg_to_check_it_4_cnu_24_in_1, msg_to_check_it_4_cnu_24_in_2, msg_to_check_it_4_cnu_24_in_3, msg_to_check_it_4_cnu_24_in_4, msg_to_check_it_4_cnu_24_in_5, msg_to_check_it_4_cnu_25_in_0, msg_to_check_it_4_cnu_25_in_1, msg_to_check_it_4_cnu_25_in_2, msg_to_check_it_4_cnu_25_in_3, msg_to_check_it_4_cnu_25_in_4, msg_to_check_it_4_cnu_25_in_5, msg_to_check_it_4_cnu_26_in_0, msg_to_check_it_4_cnu_26_in_1, msg_to_check_it_4_cnu_26_in_2, msg_to_check_it_4_cnu_26_in_3, msg_to_check_it_4_cnu_26_in_4, msg_to_check_it_4_cnu_26_in_5, msg_to_check_it_4_cnu_27_in_0, msg_to_check_it_4_cnu_27_in_1, msg_to_check_it_4_cnu_27_in_2, msg_to_check_it_4_cnu_27_in_3, msg_to_check_it_4_cnu_27_in_4, msg_to_check_it_4_cnu_27_in_5, msg_to_check_it_4_cnu_28_in_0, msg_to_check_it_4_cnu_28_in_1, msg_to_check_it_4_cnu_28_in_2, msg_to_check_it_4_cnu_28_in_3, msg_to_check_it_4_cnu_28_in_4, msg_to_check_it_4_cnu_28_in_5, msg_to_check_it_4_cnu_29_in_0, msg_to_check_it_4_cnu_29_in_1, msg_to_check_it_4_cnu_29_in_2, msg_to_check_it_4_cnu_29_in_3, msg_to_check_it_4_cnu_29_in_4, msg_to_check_it_4_cnu_29_in_5, msg_to_check_it_4_cnu_30_in_0, msg_to_check_it_4_cnu_30_in_1, msg_to_check_it_4_cnu_30_in_2, msg_to_check_it_4_cnu_30_in_3, msg_to_check_it_4_cnu_30_in_4, msg_to_check_it_4_cnu_30_in_5, msg_to_check_it_4_cnu_31_in_0, msg_to_check_it_4_cnu_31_in_1, msg_to_check_it_4_cnu_31_in_2, msg_to_check_it_4_cnu_31_in_3, msg_to_check_it_4_cnu_31_in_4, msg_to_check_it_4_cnu_31_in_5, msg_to_check_it_4_cnu_32_in_0, msg_to_check_it_4_cnu_32_in_1, msg_to_check_it_4_cnu_32_in_2, msg_to_check_it_4_cnu_32_in_3, msg_to_check_it_4_cnu_32_in_4, msg_to_check_it_4_cnu_32_in_5, msg_to_check_it_4_cnu_33_in_0, msg_to_check_it_4_cnu_33_in_1, msg_to_check_it_4_cnu_33_in_2, msg_to_check_it_4_cnu_33_in_3, msg_to_check_it_4_cnu_33_in_4, msg_to_check_it_4_cnu_33_in_5, msg_to_check_it_4_cnu_34_in_0, msg_to_check_it_4_cnu_34_in_1, msg_to_check_it_4_cnu_34_in_2, msg_to_check_it_4_cnu_34_in_3, msg_to_check_it_4_cnu_34_in_4, msg_to_check_it_4_cnu_34_in_5, msg_to_check_it_4_cnu_35_in_0, msg_to_check_it_4_cnu_35_in_1, msg_to_check_it_4_cnu_35_in_2, msg_to_check_it_4_cnu_35_in_3, msg_to_check_it_4_cnu_35_in_4, msg_to_check_it_4_cnu_35_in_5, msg_to_check_it_4_cnu_36_in_0, msg_to_check_it_4_cnu_36_in_1, msg_to_check_it_4_cnu_36_in_2, msg_to_check_it_4_cnu_36_in_3, msg_to_check_it_4_cnu_36_in_4, msg_to_check_it_4_cnu_36_in_5, msg_to_check_it_4_cnu_37_in_0, msg_to_check_it_4_cnu_37_in_1, msg_to_check_it_4_cnu_37_in_2, msg_to_check_it_4_cnu_37_in_3, msg_to_check_it_4_cnu_37_in_4, msg_to_check_it_4_cnu_37_in_5, msg_to_check_it_4_cnu_38_in_0, msg_to_check_it_4_cnu_38_in_1, msg_to_check_it_4_cnu_38_in_2, msg_to_check_it_4_cnu_38_in_3, msg_to_check_it_4_cnu_38_in_4, msg_to_check_it_4_cnu_38_in_5, msg_to_check_it_4_cnu_39_in_0, msg_to_check_it_4_cnu_39_in_1, msg_to_check_it_4_cnu_39_in_2, msg_to_check_it_4_cnu_39_in_3, msg_to_check_it_4_cnu_39_in_4, msg_to_check_it_4_cnu_39_in_5, msg_to_check_it_4_cnu_40_in_0, msg_to_check_it_4_cnu_40_in_1, msg_to_check_it_4_cnu_40_in_2, msg_to_check_it_4_cnu_40_in_3, msg_to_check_it_4_cnu_40_in_4, msg_to_check_it_4_cnu_40_in_5, msg_to_check_it_4_cnu_41_in_0, msg_to_check_it_4_cnu_41_in_1, msg_to_check_it_4_cnu_41_in_2, msg_to_check_it_4_cnu_41_in_3, msg_to_check_it_4_cnu_41_in_4, msg_to_check_it_4_cnu_41_in_5, msg_to_check_it_4_cnu_42_in_0, msg_to_check_it_4_cnu_42_in_1, msg_to_check_it_4_cnu_42_in_2, msg_to_check_it_4_cnu_42_in_3, msg_to_check_it_4_cnu_42_in_4, msg_to_check_it_4_cnu_42_in_5, msg_to_check_it_4_cnu_43_in_0, msg_to_check_it_4_cnu_43_in_1, msg_to_check_it_4_cnu_43_in_2, msg_to_check_it_4_cnu_43_in_3, msg_to_check_it_4_cnu_43_in_4, msg_to_check_it_4_cnu_43_in_5, msg_to_check_it_4_cnu_44_in_0, msg_to_check_it_4_cnu_44_in_1, msg_to_check_it_4_cnu_44_in_2, msg_to_check_it_4_cnu_44_in_3, msg_to_check_it_4_cnu_44_in_4, msg_to_check_it_4_cnu_44_in_5, msg_to_check_it_4_cnu_45_in_0, msg_to_check_it_4_cnu_45_in_1, msg_to_check_it_4_cnu_45_in_2, msg_to_check_it_4_cnu_45_in_3, msg_to_check_it_4_cnu_45_in_4, msg_to_check_it_4_cnu_45_in_5, msg_to_check_it_4_cnu_46_in_0, msg_to_check_it_4_cnu_46_in_1, msg_to_check_it_4_cnu_46_in_2, msg_to_check_it_4_cnu_46_in_3, msg_to_check_it_4_cnu_46_in_4, msg_to_check_it_4_cnu_46_in_5, msg_to_check_it_4_cnu_47_in_0, msg_to_check_it_4_cnu_47_in_1, msg_to_check_it_4_cnu_47_in_2, msg_to_check_it_4_cnu_47_in_3, msg_to_check_it_4_cnu_47_in_4, msg_to_check_it_4_cnu_47_in_5, msg_to_check_it_4_cnu_48_in_0, msg_to_check_it_4_cnu_48_in_1, msg_to_check_it_4_cnu_48_in_2, msg_to_check_it_4_cnu_48_in_3, msg_to_check_it_4_cnu_48_in_4, msg_to_check_it_4_cnu_48_in_5, msg_to_check_it_4_cnu_49_in_0, msg_to_check_it_4_cnu_49_in_1, msg_to_check_it_4_cnu_49_in_2, msg_to_check_it_4_cnu_49_in_3, msg_to_check_it_4_cnu_49_in_4, msg_to_check_it_4_cnu_49_in_5, msg_to_check_it_4_cnu_50_in_0, msg_to_check_it_4_cnu_50_in_1, msg_to_check_it_4_cnu_50_in_2, msg_to_check_it_4_cnu_50_in_3, msg_to_check_it_4_cnu_50_in_4, msg_to_check_it_4_cnu_50_in_5, msg_to_check_it_4_cnu_51_in_0, msg_to_check_it_4_cnu_51_in_1, msg_to_check_it_4_cnu_51_in_2, msg_to_check_it_4_cnu_51_in_3, msg_to_check_it_4_cnu_51_in_4, msg_to_check_it_4_cnu_51_in_5, msg_to_check_it_4_cnu_52_in_0, msg_to_check_it_4_cnu_52_in_1, msg_to_check_it_4_cnu_52_in_2, msg_to_check_it_4_cnu_52_in_3, msg_to_check_it_4_cnu_52_in_4, msg_to_check_it_4_cnu_52_in_5, msg_to_check_it_4_cnu_53_in_0, msg_to_check_it_4_cnu_53_in_1, msg_to_check_it_4_cnu_53_in_2, msg_to_check_it_4_cnu_53_in_3, msg_to_check_it_4_cnu_53_in_4, msg_to_check_it_4_cnu_53_in_5, msg_to_check_it_4_cnu_54_in_0, msg_to_check_it_4_cnu_54_in_1, msg_to_check_it_4_cnu_54_in_2, msg_to_check_it_4_cnu_54_in_3, msg_to_check_it_4_cnu_54_in_4, msg_to_check_it_4_cnu_54_in_5, msg_to_check_it_4_cnu_55_in_0, msg_to_check_it_4_cnu_55_in_1, msg_to_check_it_4_cnu_55_in_2, msg_to_check_it_4_cnu_55_in_3, msg_to_check_it_4_cnu_55_in_4, msg_to_check_it_4_cnu_55_in_5, msg_to_check_it_4_cnu_56_in_0, msg_to_check_it_4_cnu_56_in_1, msg_to_check_it_4_cnu_56_in_2, msg_to_check_it_4_cnu_56_in_3, msg_to_check_it_4_cnu_56_in_4, msg_to_check_it_4_cnu_56_in_5, msg_to_check_it_4_cnu_57_in_0, msg_to_check_it_4_cnu_57_in_1, msg_to_check_it_4_cnu_57_in_2, msg_to_check_it_4_cnu_57_in_3, msg_to_check_it_4_cnu_57_in_4, msg_to_check_it_4_cnu_57_in_5, msg_to_check_it_4_cnu_58_in_0, msg_to_check_it_4_cnu_58_in_1, msg_to_check_it_4_cnu_58_in_2, msg_to_check_it_4_cnu_58_in_3, msg_to_check_it_4_cnu_58_in_4, msg_to_check_it_4_cnu_58_in_5, msg_to_check_it_4_cnu_59_in_0, msg_to_check_it_4_cnu_59_in_1, msg_to_check_it_4_cnu_59_in_2, msg_to_check_it_4_cnu_59_in_3, msg_to_check_it_4_cnu_59_in_4, msg_to_check_it_4_cnu_59_in_5, msg_to_check_it_4_cnu_60_in_0, msg_to_check_it_4_cnu_60_in_1, msg_to_check_it_4_cnu_60_in_2, msg_to_check_it_4_cnu_60_in_3, msg_to_check_it_4_cnu_60_in_4, msg_to_check_it_4_cnu_60_in_5, msg_to_check_it_4_cnu_61_in_0, msg_to_check_it_4_cnu_61_in_1, msg_to_check_it_4_cnu_61_in_2, msg_to_check_it_4_cnu_61_in_3, msg_to_check_it_4_cnu_61_in_4, msg_to_check_it_4_cnu_61_in_5, msg_to_check_it_4_cnu_62_in_0, msg_to_check_it_4_cnu_62_in_1, msg_to_check_it_4_cnu_62_in_2, msg_to_check_it_4_cnu_62_in_3, msg_to_check_it_4_cnu_62_in_4, msg_to_check_it_4_cnu_62_in_5, msg_to_check_it_4_cnu_63_in_0, msg_to_check_it_4_cnu_63_in_1, msg_to_check_it_4_cnu_63_in_2, msg_to_check_it_4_cnu_63_in_3, msg_to_check_it_4_cnu_63_in_4, msg_to_check_it_4_cnu_63_in_5, msg_to_check_it_4_cnu_64_in_0, msg_to_check_it_4_cnu_64_in_1, msg_to_check_it_4_cnu_64_in_2, msg_to_check_it_4_cnu_64_in_3, msg_to_check_it_4_cnu_64_in_4, msg_to_check_it_4_cnu_64_in_5, msg_to_check_it_4_cnu_65_in_0, msg_to_check_it_4_cnu_65_in_1, msg_to_check_it_4_cnu_65_in_2, msg_to_check_it_4_cnu_65_in_3, msg_to_check_it_4_cnu_65_in_4, msg_to_check_it_4_cnu_65_in_5, msg_to_check_it_4_cnu_66_in_0, msg_to_check_it_4_cnu_66_in_1, msg_to_check_it_4_cnu_66_in_2, msg_to_check_it_4_cnu_66_in_3, msg_to_check_it_4_cnu_66_in_4, msg_to_check_it_4_cnu_66_in_5, msg_to_check_it_4_cnu_67_in_0, msg_to_check_it_4_cnu_67_in_1, msg_to_check_it_4_cnu_67_in_2, msg_to_check_it_4_cnu_67_in_3, msg_to_check_it_4_cnu_67_in_4, msg_to_check_it_4_cnu_67_in_5, msg_to_check_it_4_cnu_68_in_0, msg_to_check_it_4_cnu_68_in_1, msg_to_check_it_4_cnu_68_in_2, msg_to_check_it_4_cnu_68_in_3, msg_to_check_it_4_cnu_68_in_4, msg_to_check_it_4_cnu_68_in_5, msg_to_check_it_4_cnu_69_in_0, msg_to_check_it_4_cnu_69_in_1, msg_to_check_it_4_cnu_69_in_2, msg_to_check_it_4_cnu_69_in_3, msg_to_check_it_4_cnu_69_in_4, msg_to_check_it_4_cnu_69_in_5, msg_to_check_it_4_cnu_70_in_0, msg_to_check_it_4_cnu_70_in_1, msg_to_check_it_4_cnu_70_in_2, msg_to_check_it_4_cnu_70_in_3, msg_to_check_it_4_cnu_70_in_4, msg_to_check_it_4_cnu_70_in_5, msg_to_check_it_4_cnu_71_in_0, msg_to_check_it_4_cnu_71_in_1, msg_to_check_it_4_cnu_71_in_2, msg_to_check_it_4_cnu_71_in_3, msg_to_check_it_4_cnu_71_in_4, msg_to_check_it_4_cnu_71_in_5, msg_to_check_it_4_cnu_72_in_0, msg_to_check_it_4_cnu_72_in_1, msg_to_check_it_4_cnu_72_in_2, msg_to_check_it_4_cnu_72_in_3, msg_to_check_it_4_cnu_72_in_4, msg_to_check_it_4_cnu_72_in_5, msg_to_check_it_4_cnu_73_in_0, msg_to_check_it_4_cnu_73_in_1, msg_to_check_it_4_cnu_73_in_2, msg_to_check_it_4_cnu_73_in_3, msg_to_check_it_4_cnu_73_in_4, msg_to_check_it_4_cnu_73_in_5, msg_to_check_it_4_cnu_74_in_0, msg_to_check_it_4_cnu_74_in_1, msg_to_check_it_4_cnu_74_in_2, msg_to_check_it_4_cnu_74_in_3, msg_to_check_it_4_cnu_74_in_4, msg_to_check_it_4_cnu_74_in_5, msg_to_check_it_4_cnu_75_in_0, msg_to_check_it_4_cnu_75_in_1, msg_to_check_it_4_cnu_75_in_2, msg_to_check_it_4_cnu_75_in_3, msg_to_check_it_4_cnu_75_in_4, msg_to_check_it_4_cnu_75_in_5, msg_to_check_it_4_cnu_76_in_0, msg_to_check_it_4_cnu_76_in_1, msg_to_check_it_4_cnu_76_in_2, msg_to_check_it_4_cnu_76_in_3, msg_to_check_it_4_cnu_76_in_4, msg_to_check_it_4_cnu_76_in_5, msg_to_check_it_4_cnu_77_in_0, msg_to_check_it_4_cnu_77_in_1, msg_to_check_it_4_cnu_77_in_2, msg_to_check_it_4_cnu_77_in_3, msg_to_check_it_4_cnu_77_in_4, msg_to_check_it_4_cnu_77_in_5, msg_to_check_it_4_cnu_78_in_0, msg_to_check_it_4_cnu_78_in_1, msg_to_check_it_4_cnu_78_in_2, msg_to_check_it_4_cnu_78_in_3, msg_to_check_it_4_cnu_78_in_4, msg_to_check_it_4_cnu_78_in_5, msg_to_check_it_4_cnu_79_in_0, msg_to_check_it_4_cnu_79_in_1, msg_to_check_it_4_cnu_79_in_2, msg_to_check_it_4_cnu_79_in_3, msg_to_check_it_4_cnu_79_in_4, msg_to_check_it_4_cnu_79_in_5, msg_to_check_it_4_cnu_80_in_0, msg_to_check_it_4_cnu_80_in_1, msg_to_check_it_4_cnu_80_in_2, msg_to_check_it_4_cnu_80_in_3, msg_to_check_it_4_cnu_80_in_4, msg_to_check_it_4_cnu_80_in_5, msg_to_check_it_4_cnu_81_in_0, msg_to_check_it_4_cnu_81_in_1, msg_to_check_it_4_cnu_81_in_2, msg_to_check_it_4_cnu_81_in_3, msg_to_check_it_4_cnu_81_in_4, msg_to_check_it_4_cnu_81_in_5, msg_to_check_it_4_cnu_82_in_0, msg_to_check_it_4_cnu_82_in_1, msg_to_check_it_4_cnu_82_in_2, msg_to_check_it_4_cnu_82_in_3, msg_to_check_it_4_cnu_82_in_4, msg_to_check_it_4_cnu_82_in_5, msg_to_check_it_4_cnu_83_in_0, msg_to_check_it_4_cnu_83_in_1, msg_to_check_it_4_cnu_83_in_2, msg_to_check_it_4_cnu_83_in_3, msg_to_check_it_4_cnu_83_in_4, msg_to_check_it_4_cnu_83_in_5, msg_to_check_it_4_cnu_84_in_0, msg_to_check_it_4_cnu_84_in_1, msg_to_check_it_4_cnu_84_in_2, msg_to_check_it_4_cnu_84_in_3, msg_to_check_it_4_cnu_84_in_4, msg_to_check_it_4_cnu_84_in_5, msg_to_check_it_4_cnu_85_in_0, msg_to_check_it_4_cnu_85_in_1, msg_to_check_it_4_cnu_85_in_2, msg_to_check_it_4_cnu_85_in_3, msg_to_check_it_4_cnu_85_in_4, msg_to_check_it_4_cnu_85_in_5, msg_to_check_it_4_cnu_86_in_0, msg_to_check_it_4_cnu_86_in_1, msg_to_check_it_4_cnu_86_in_2, msg_to_check_it_4_cnu_86_in_3, msg_to_check_it_4_cnu_86_in_4, msg_to_check_it_4_cnu_86_in_5, msg_to_check_it_4_cnu_87_in_0, msg_to_check_it_4_cnu_87_in_1, msg_to_check_it_4_cnu_87_in_2, msg_to_check_it_4_cnu_87_in_3, msg_to_check_it_4_cnu_87_in_4, msg_to_check_it_4_cnu_87_in_5, msg_to_check_it_4_cnu_88_in_0, msg_to_check_it_4_cnu_88_in_1, msg_to_check_it_4_cnu_88_in_2, msg_to_check_it_4_cnu_88_in_3, msg_to_check_it_4_cnu_88_in_4, msg_to_check_it_4_cnu_88_in_5, msg_to_check_it_4_cnu_89_in_0, msg_to_check_it_4_cnu_89_in_1, msg_to_check_it_4_cnu_89_in_2, msg_to_check_it_4_cnu_89_in_3, msg_to_check_it_4_cnu_89_in_4, msg_to_check_it_4_cnu_89_in_5, msg_to_check_it_4_cnu_90_in_0, msg_to_check_it_4_cnu_90_in_1, msg_to_check_it_4_cnu_90_in_2, msg_to_check_it_4_cnu_90_in_3, msg_to_check_it_4_cnu_90_in_4, msg_to_check_it_4_cnu_90_in_5, msg_to_check_it_4_cnu_91_in_0, msg_to_check_it_4_cnu_91_in_1, msg_to_check_it_4_cnu_91_in_2, msg_to_check_it_4_cnu_91_in_3, msg_to_check_it_4_cnu_91_in_4, msg_to_check_it_4_cnu_91_in_5, msg_to_check_it_4_cnu_92_in_0, msg_to_check_it_4_cnu_92_in_1, msg_to_check_it_4_cnu_92_in_2, msg_to_check_it_4_cnu_92_in_3, msg_to_check_it_4_cnu_92_in_4, msg_to_check_it_4_cnu_92_in_5, msg_to_check_it_4_cnu_93_in_0, msg_to_check_it_4_cnu_93_in_1, msg_to_check_it_4_cnu_93_in_2, msg_to_check_it_4_cnu_93_in_3, msg_to_check_it_4_cnu_93_in_4, msg_to_check_it_4_cnu_93_in_5, msg_to_check_it_4_cnu_94_in_0, msg_to_check_it_4_cnu_94_in_1, msg_to_check_it_4_cnu_94_in_2, msg_to_check_it_4_cnu_94_in_3, msg_to_check_it_4_cnu_94_in_4, msg_to_check_it_4_cnu_94_in_5, msg_to_check_it_4_cnu_95_in_0, msg_to_check_it_4_cnu_95_in_1, msg_to_check_it_4_cnu_95_in_2, msg_to_check_it_4_cnu_95_in_3, msg_to_check_it_4_cnu_95_in_4, msg_to_check_it_4_cnu_95_in_5, msg_to_check_it_4_cnu_96_in_0, msg_to_check_it_4_cnu_96_in_1, msg_to_check_it_4_cnu_96_in_2, msg_to_check_it_4_cnu_96_in_3, msg_to_check_it_4_cnu_96_in_4, msg_to_check_it_4_cnu_96_in_5, msg_to_check_it_4_cnu_97_in_0, msg_to_check_it_4_cnu_97_in_1, msg_to_check_it_4_cnu_97_in_2, msg_to_check_it_4_cnu_97_in_3, msg_to_check_it_4_cnu_97_in_4, msg_to_check_it_4_cnu_97_in_5, msg_to_check_it_4_cnu_98_in_0, msg_to_check_it_4_cnu_98_in_1, msg_to_check_it_4_cnu_98_in_2, msg_to_check_it_4_cnu_98_in_3, msg_to_check_it_4_cnu_98_in_4, msg_to_check_it_4_cnu_98_in_5, msg_to_check_it_5_cnu_0_in_0, msg_to_check_it_5_cnu_0_in_1, msg_to_check_it_5_cnu_0_in_2, msg_to_check_it_5_cnu_0_in_3, msg_to_check_it_5_cnu_0_in_4, msg_to_check_it_5_cnu_0_in_5, msg_to_check_it_5_cnu_1_in_0, msg_to_check_it_5_cnu_1_in_1, msg_to_check_it_5_cnu_1_in_2, msg_to_check_it_5_cnu_1_in_3, msg_to_check_it_5_cnu_1_in_4, msg_to_check_it_5_cnu_1_in_5, msg_to_check_it_5_cnu_2_in_0, msg_to_check_it_5_cnu_2_in_1, msg_to_check_it_5_cnu_2_in_2, msg_to_check_it_5_cnu_2_in_3, msg_to_check_it_5_cnu_2_in_4, msg_to_check_it_5_cnu_2_in_5, msg_to_check_it_5_cnu_3_in_0, msg_to_check_it_5_cnu_3_in_1, msg_to_check_it_5_cnu_3_in_2, msg_to_check_it_5_cnu_3_in_3, msg_to_check_it_5_cnu_3_in_4, msg_to_check_it_5_cnu_3_in_5, msg_to_check_it_5_cnu_4_in_0, msg_to_check_it_5_cnu_4_in_1, msg_to_check_it_5_cnu_4_in_2, msg_to_check_it_5_cnu_4_in_3, msg_to_check_it_5_cnu_4_in_4, msg_to_check_it_5_cnu_4_in_5, msg_to_check_it_5_cnu_5_in_0, msg_to_check_it_5_cnu_5_in_1, msg_to_check_it_5_cnu_5_in_2, msg_to_check_it_5_cnu_5_in_3, msg_to_check_it_5_cnu_5_in_4, msg_to_check_it_5_cnu_5_in_5, msg_to_check_it_5_cnu_6_in_0, msg_to_check_it_5_cnu_6_in_1, msg_to_check_it_5_cnu_6_in_2, msg_to_check_it_5_cnu_6_in_3, msg_to_check_it_5_cnu_6_in_4, msg_to_check_it_5_cnu_6_in_5, msg_to_check_it_5_cnu_7_in_0, msg_to_check_it_5_cnu_7_in_1, msg_to_check_it_5_cnu_7_in_2, msg_to_check_it_5_cnu_7_in_3, msg_to_check_it_5_cnu_7_in_4, msg_to_check_it_5_cnu_7_in_5, msg_to_check_it_5_cnu_8_in_0, msg_to_check_it_5_cnu_8_in_1, msg_to_check_it_5_cnu_8_in_2, msg_to_check_it_5_cnu_8_in_3, msg_to_check_it_5_cnu_8_in_4, msg_to_check_it_5_cnu_8_in_5, msg_to_check_it_5_cnu_9_in_0, msg_to_check_it_5_cnu_9_in_1, msg_to_check_it_5_cnu_9_in_2, msg_to_check_it_5_cnu_9_in_3, msg_to_check_it_5_cnu_9_in_4, msg_to_check_it_5_cnu_9_in_5, msg_to_check_it_5_cnu_10_in_0, msg_to_check_it_5_cnu_10_in_1, msg_to_check_it_5_cnu_10_in_2, msg_to_check_it_5_cnu_10_in_3, msg_to_check_it_5_cnu_10_in_4, msg_to_check_it_5_cnu_10_in_5, msg_to_check_it_5_cnu_11_in_0, msg_to_check_it_5_cnu_11_in_1, msg_to_check_it_5_cnu_11_in_2, msg_to_check_it_5_cnu_11_in_3, msg_to_check_it_5_cnu_11_in_4, msg_to_check_it_5_cnu_11_in_5, msg_to_check_it_5_cnu_12_in_0, msg_to_check_it_5_cnu_12_in_1, msg_to_check_it_5_cnu_12_in_2, msg_to_check_it_5_cnu_12_in_3, msg_to_check_it_5_cnu_12_in_4, msg_to_check_it_5_cnu_12_in_5, msg_to_check_it_5_cnu_13_in_0, msg_to_check_it_5_cnu_13_in_1, msg_to_check_it_5_cnu_13_in_2, msg_to_check_it_5_cnu_13_in_3, msg_to_check_it_5_cnu_13_in_4, msg_to_check_it_5_cnu_13_in_5, msg_to_check_it_5_cnu_14_in_0, msg_to_check_it_5_cnu_14_in_1, msg_to_check_it_5_cnu_14_in_2, msg_to_check_it_5_cnu_14_in_3, msg_to_check_it_5_cnu_14_in_4, msg_to_check_it_5_cnu_14_in_5, msg_to_check_it_5_cnu_15_in_0, msg_to_check_it_5_cnu_15_in_1, msg_to_check_it_5_cnu_15_in_2, msg_to_check_it_5_cnu_15_in_3, msg_to_check_it_5_cnu_15_in_4, msg_to_check_it_5_cnu_15_in_5, msg_to_check_it_5_cnu_16_in_0, msg_to_check_it_5_cnu_16_in_1, msg_to_check_it_5_cnu_16_in_2, msg_to_check_it_5_cnu_16_in_3, msg_to_check_it_5_cnu_16_in_4, msg_to_check_it_5_cnu_16_in_5, msg_to_check_it_5_cnu_17_in_0, msg_to_check_it_5_cnu_17_in_1, msg_to_check_it_5_cnu_17_in_2, msg_to_check_it_5_cnu_17_in_3, msg_to_check_it_5_cnu_17_in_4, msg_to_check_it_5_cnu_17_in_5, msg_to_check_it_5_cnu_18_in_0, msg_to_check_it_5_cnu_18_in_1, msg_to_check_it_5_cnu_18_in_2, msg_to_check_it_5_cnu_18_in_3, msg_to_check_it_5_cnu_18_in_4, msg_to_check_it_5_cnu_18_in_5, msg_to_check_it_5_cnu_19_in_0, msg_to_check_it_5_cnu_19_in_1, msg_to_check_it_5_cnu_19_in_2, msg_to_check_it_5_cnu_19_in_3, msg_to_check_it_5_cnu_19_in_4, msg_to_check_it_5_cnu_19_in_5, msg_to_check_it_5_cnu_20_in_0, msg_to_check_it_5_cnu_20_in_1, msg_to_check_it_5_cnu_20_in_2, msg_to_check_it_5_cnu_20_in_3, msg_to_check_it_5_cnu_20_in_4, msg_to_check_it_5_cnu_20_in_5, msg_to_check_it_5_cnu_21_in_0, msg_to_check_it_5_cnu_21_in_1, msg_to_check_it_5_cnu_21_in_2, msg_to_check_it_5_cnu_21_in_3, msg_to_check_it_5_cnu_21_in_4, msg_to_check_it_5_cnu_21_in_5, msg_to_check_it_5_cnu_22_in_0, msg_to_check_it_5_cnu_22_in_1, msg_to_check_it_5_cnu_22_in_2, msg_to_check_it_5_cnu_22_in_3, msg_to_check_it_5_cnu_22_in_4, msg_to_check_it_5_cnu_22_in_5, msg_to_check_it_5_cnu_23_in_0, msg_to_check_it_5_cnu_23_in_1, msg_to_check_it_5_cnu_23_in_2, msg_to_check_it_5_cnu_23_in_3, msg_to_check_it_5_cnu_23_in_4, msg_to_check_it_5_cnu_23_in_5, msg_to_check_it_5_cnu_24_in_0, msg_to_check_it_5_cnu_24_in_1, msg_to_check_it_5_cnu_24_in_2, msg_to_check_it_5_cnu_24_in_3, msg_to_check_it_5_cnu_24_in_4, msg_to_check_it_5_cnu_24_in_5, msg_to_check_it_5_cnu_25_in_0, msg_to_check_it_5_cnu_25_in_1, msg_to_check_it_5_cnu_25_in_2, msg_to_check_it_5_cnu_25_in_3, msg_to_check_it_5_cnu_25_in_4, msg_to_check_it_5_cnu_25_in_5, msg_to_check_it_5_cnu_26_in_0, msg_to_check_it_5_cnu_26_in_1, msg_to_check_it_5_cnu_26_in_2, msg_to_check_it_5_cnu_26_in_3, msg_to_check_it_5_cnu_26_in_4, msg_to_check_it_5_cnu_26_in_5, msg_to_check_it_5_cnu_27_in_0, msg_to_check_it_5_cnu_27_in_1, msg_to_check_it_5_cnu_27_in_2, msg_to_check_it_5_cnu_27_in_3, msg_to_check_it_5_cnu_27_in_4, msg_to_check_it_5_cnu_27_in_5, msg_to_check_it_5_cnu_28_in_0, msg_to_check_it_5_cnu_28_in_1, msg_to_check_it_5_cnu_28_in_2, msg_to_check_it_5_cnu_28_in_3, msg_to_check_it_5_cnu_28_in_4, msg_to_check_it_5_cnu_28_in_5, msg_to_check_it_5_cnu_29_in_0, msg_to_check_it_5_cnu_29_in_1, msg_to_check_it_5_cnu_29_in_2, msg_to_check_it_5_cnu_29_in_3, msg_to_check_it_5_cnu_29_in_4, msg_to_check_it_5_cnu_29_in_5, msg_to_check_it_5_cnu_30_in_0, msg_to_check_it_5_cnu_30_in_1, msg_to_check_it_5_cnu_30_in_2, msg_to_check_it_5_cnu_30_in_3, msg_to_check_it_5_cnu_30_in_4, msg_to_check_it_5_cnu_30_in_5, msg_to_check_it_5_cnu_31_in_0, msg_to_check_it_5_cnu_31_in_1, msg_to_check_it_5_cnu_31_in_2, msg_to_check_it_5_cnu_31_in_3, msg_to_check_it_5_cnu_31_in_4, msg_to_check_it_5_cnu_31_in_5, msg_to_check_it_5_cnu_32_in_0, msg_to_check_it_5_cnu_32_in_1, msg_to_check_it_5_cnu_32_in_2, msg_to_check_it_5_cnu_32_in_3, msg_to_check_it_5_cnu_32_in_4, msg_to_check_it_5_cnu_32_in_5, msg_to_check_it_5_cnu_33_in_0, msg_to_check_it_5_cnu_33_in_1, msg_to_check_it_5_cnu_33_in_2, msg_to_check_it_5_cnu_33_in_3, msg_to_check_it_5_cnu_33_in_4, msg_to_check_it_5_cnu_33_in_5, msg_to_check_it_5_cnu_34_in_0, msg_to_check_it_5_cnu_34_in_1, msg_to_check_it_5_cnu_34_in_2, msg_to_check_it_5_cnu_34_in_3, msg_to_check_it_5_cnu_34_in_4, msg_to_check_it_5_cnu_34_in_5, msg_to_check_it_5_cnu_35_in_0, msg_to_check_it_5_cnu_35_in_1, msg_to_check_it_5_cnu_35_in_2, msg_to_check_it_5_cnu_35_in_3, msg_to_check_it_5_cnu_35_in_4, msg_to_check_it_5_cnu_35_in_5, msg_to_check_it_5_cnu_36_in_0, msg_to_check_it_5_cnu_36_in_1, msg_to_check_it_5_cnu_36_in_2, msg_to_check_it_5_cnu_36_in_3, msg_to_check_it_5_cnu_36_in_4, msg_to_check_it_5_cnu_36_in_5, msg_to_check_it_5_cnu_37_in_0, msg_to_check_it_5_cnu_37_in_1, msg_to_check_it_5_cnu_37_in_2, msg_to_check_it_5_cnu_37_in_3, msg_to_check_it_5_cnu_37_in_4, msg_to_check_it_5_cnu_37_in_5, msg_to_check_it_5_cnu_38_in_0, msg_to_check_it_5_cnu_38_in_1, msg_to_check_it_5_cnu_38_in_2, msg_to_check_it_5_cnu_38_in_3, msg_to_check_it_5_cnu_38_in_4, msg_to_check_it_5_cnu_38_in_5, msg_to_check_it_5_cnu_39_in_0, msg_to_check_it_5_cnu_39_in_1, msg_to_check_it_5_cnu_39_in_2, msg_to_check_it_5_cnu_39_in_3, msg_to_check_it_5_cnu_39_in_4, msg_to_check_it_5_cnu_39_in_5, msg_to_check_it_5_cnu_40_in_0, msg_to_check_it_5_cnu_40_in_1, msg_to_check_it_5_cnu_40_in_2, msg_to_check_it_5_cnu_40_in_3, msg_to_check_it_5_cnu_40_in_4, msg_to_check_it_5_cnu_40_in_5, msg_to_check_it_5_cnu_41_in_0, msg_to_check_it_5_cnu_41_in_1, msg_to_check_it_5_cnu_41_in_2, msg_to_check_it_5_cnu_41_in_3, msg_to_check_it_5_cnu_41_in_4, msg_to_check_it_5_cnu_41_in_5, msg_to_check_it_5_cnu_42_in_0, msg_to_check_it_5_cnu_42_in_1, msg_to_check_it_5_cnu_42_in_2, msg_to_check_it_5_cnu_42_in_3, msg_to_check_it_5_cnu_42_in_4, msg_to_check_it_5_cnu_42_in_5, msg_to_check_it_5_cnu_43_in_0, msg_to_check_it_5_cnu_43_in_1, msg_to_check_it_5_cnu_43_in_2, msg_to_check_it_5_cnu_43_in_3, msg_to_check_it_5_cnu_43_in_4, msg_to_check_it_5_cnu_43_in_5, msg_to_check_it_5_cnu_44_in_0, msg_to_check_it_5_cnu_44_in_1, msg_to_check_it_5_cnu_44_in_2, msg_to_check_it_5_cnu_44_in_3, msg_to_check_it_5_cnu_44_in_4, msg_to_check_it_5_cnu_44_in_5, msg_to_check_it_5_cnu_45_in_0, msg_to_check_it_5_cnu_45_in_1, msg_to_check_it_5_cnu_45_in_2, msg_to_check_it_5_cnu_45_in_3, msg_to_check_it_5_cnu_45_in_4, msg_to_check_it_5_cnu_45_in_5, msg_to_check_it_5_cnu_46_in_0, msg_to_check_it_5_cnu_46_in_1, msg_to_check_it_5_cnu_46_in_2, msg_to_check_it_5_cnu_46_in_3, msg_to_check_it_5_cnu_46_in_4, msg_to_check_it_5_cnu_46_in_5, msg_to_check_it_5_cnu_47_in_0, msg_to_check_it_5_cnu_47_in_1, msg_to_check_it_5_cnu_47_in_2, msg_to_check_it_5_cnu_47_in_3, msg_to_check_it_5_cnu_47_in_4, msg_to_check_it_5_cnu_47_in_5, msg_to_check_it_5_cnu_48_in_0, msg_to_check_it_5_cnu_48_in_1, msg_to_check_it_5_cnu_48_in_2, msg_to_check_it_5_cnu_48_in_3, msg_to_check_it_5_cnu_48_in_4, msg_to_check_it_5_cnu_48_in_5, msg_to_check_it_5_cnu_49_in_0, msg_to_check_it_5_cnu_49_in_1, msg_to_check_it_5_cnu_49_in_2, msg_to_check_it_5_cnu_49_in_3, msg_to_check_it_5_cnu_49_in_4, msg_to_check_it_5_cnu_49_in_5, msg_to_check_it_5_cnu_50_in_0, msg_to_check_it_5_cnu_50_in_1, msg_to_check_it_5_cnu_50_in_2, msg_to_check_it_5_cnu_50_in_3, msg_to_check_it_5_cnu_50_in_4, msg_to_check_it_5_cnu_50_in_5, msg_to_check_it_5_cnu_51_in_0, msg_to_check_it_5_cnu_51_in_1, msg_to_check_it_5_cnu_51_in_2, msg_to_check_it_5_cnu_51_in_3, msg_to_check_it_5_cnu_51_in_4, msg_to_check_it_5_cnu_51_in_5, msg_to_check_it_5_cnu_52_in_0, msg_to_check_it_5_cnu_52_in_1, msg_to_check_it_5_cnu_52_in_2, msg_to_check_it_5_cnu_52_in_3, msg_to_check_it_5_cnu_52_in_4, msg_to_check_it_5_cnu_52_in_5, msg_to_check_it_5_cnu_53_in_0, msg_to_check_it_5_cnu_53_in_1, msg_to_check_it_5_cnu_53_in_2, msg_to_check_it_5_cnu_53_in_3, msg_to_check_it_5_cnu_53_in_4, msg_to_check_it_5_cnu_53_in_5, msg_to_check_it_5_cnu_54_in_0, msg_to_check_it_5_cnu_54_in_1, msg_to_check_it_5_cnu_54_in_2, msg_to_check_it_5_cnu_54_in_3, msg_to_check_it_5_cnu_54_in_4, msg_to_check_it_5_cnu_54_in_5, msg_to_check_it_5_cnu_55_in_0, msg_to_check_it_5_cnu_55_in_1, msg_to_check_it_5_cnu_55_in_2, msg_to_check_it_5_cnu_55_in_3, msg_to_check_it_5_cnu_55_in_4, msg_to_check_it_5_cnu_55_in_5, msg_to_check_it_5_cnu_56_in_0, msg_to_check_it_5_cnu_56_in_1, msg_to_check_it_5_cnu_56_in_2, msg_to_check_it_5_cnu_56_in_3, msg_to_check_it_5_cnu_56_in_4, msg_to_check_it_5_cnu_56_in_5, msg_to_check_it_5_cnu_57_in_0, msg_to_check_it_5_cnu_57_in_1, msg_to_check_it_5_cnu_57_in_2, msg_to_check_it_5_cnu_57_in_3, msg_to_check_it_5_cnu_57_in_4, msg_to_check_it_5_cnu_57_in_5, msg_to_check_it_5_cnu_58_in_0, msg_to_check_it_5_cnu_58_in_1, msg_to_check_it_5_cnu_58_in_2, msg_to_check_it_5_cnu_58_in_3, msg_to_check_it_5_cnu_58_in_4, msg_to_check_it_5_cnu_58_in_5, msg_to_check_it_5_cnu_59_in_0, msg_to_check_it_5_cnu_59_in_1, msg_to_check_it_5_cnu_59_in_2, msg_to_check_it_5_cnu_59_in_3, msg_to_check_it_5_cnu_59_in_4, msg_to_check_it_5_cnu_59_in_5, msg_to_check_it_5_cnu_60_in_0, msg_to_check_it_5_cnu_60_in_1, msg_to_check_it_5_cnu_60_in_2, msg_to_check_it_5_cnu_60_in_3, msg_to_check_it_5_cnu_60_in_4, msg_to_check_it_5_cnu_60_in_5, msg_to_check_it_5_cnu_61_in_0, msg_to_check_it_5_cnu_61_in_1, msg_to_check_it_5_cnu_61_in_2, msg_to_check_it_5_cnu_61_in_3, msg_to_check_it_5_cnu_61_in_4, msg_to_check_it_5_cnu_61_in_5, msg_to_check_it_5_cnu_62_in_0, msg_to_check_it_5_cnu_62_in_1, msg_to_check_it_5_cnu_62_in_2, msg_to_check_it_5_cnu_62_in_3, msg_to_check_it_5_cnu_62_in_4, msg_to_check_it_5_cnu_62_in_5, msg_to_check_it_5_cnu_63_in_0, msg_to_check_it_5_cnu_63_in_1, msg_to_check_it_5_cnu_63_in_2, msg_to_check_it_5_cnu_63_in_3, msg_to_check_it_5_cnu_63_in_4, msg_to_check_it_5_cnu_63_in_5, msg_to_check_it_5_cnu_64_in_0, msg_to_check_it_5_cnu_64_in_1, msg_to_check_it_5_cnu_64_in_2, msg_to_check_it_5_cnu_64_in_3, msg_to_check_it_5_cnu_64_in_4, msg_to_check_it_5_cnu_64_in_5, msg_to_check_it_5_cnu_65_in_0, msg_to_check_it_5_cnu_65_in_1, msg_to_check_it_5_cnu_65_in_2, msg_to_check_it_5_cnu_65_in_3, msg_to_check_it_5_cnu_65_in_4, msg_to_check_it_5_cnu_65_in_5, msg_to_check_it_5_cnu_66_in_0, msg_to_check_it_5_cnu_66_in_1, msg_to_check_it_5_cnu_66_in_2, msg_to_check_it_5_cnu_66_in_3, msg_to_check_it_5_cnu_66_in_4, msg_to_check_it_5_cnu_66_in_5, msg_to_check_it_5_cnu_67_in_0, msg_to_check_it_5_cnu_67_in_1, msg_to_check_it_5_cnu_67_in_2, msg_to_check_it_5_cnu_67_in_3, msg_to_check_it_5_cnu_67_in_4, msg_to_check_it_5_cnu_67_in_5, msg_to_check_it_5_cnu_68_in_0, msg_to_check_it_5_cnu_68_in_1, msg_to_check_it_5_cnu_68_in_2, msg_to_check_it_5_cnu_68_in_3, msg_to_check_it_5_cnu_68_in_4, msg_to_check_it_5_cnu_68_in_5, msg_to_check_it_5_cnu_69_in_0, msg_to_check_it_5_cnu_69_in_1, msg_to_check_it_5_cnu_69_in_2, msg_to_check_it_5_cnu_69_in_3, msg_to_check_it_5_cnu_69_in_4, msg_to_check_it_5_cnu_69_in_5, msg_to_check_it_5_cnu_70_in_0, msg_to_check_it_5_cnu_70_in_1, msg_to_check_it_5_cnu_70_in_2, msg_to_check_it_5_cnu_70_in_3, msg_to_check_it_5_cnu_70_in_4, msg_to_check_it_5_cnu_70_in_5, msg_to_check_it_5_cnu_71_in_0, msg_to_check_it_5_cnu_71_in_1, msg_to_check_it_5_cnu_71_in_2, msg_to_check_it_5_cnu_71_in_3, msg_to_check_it_5_cnu_71_in_4, msg_to_check_it_5_cnu_71_in_5, msg_to_check_it_5_cnu_72_in_0, msg_to_check_it_5_cnu_72_in_1, msg_to_check_it_5_cnu_72_in_2, msg_to_check_it_5_cnu_72_in_3, msg_to_check_it_5_cnu_72_in_4, msg_to_check_it_5_cnu_72_in_5, msg_to_check_it_5_cnu_73_in_0, msg_to_check_it_5_cnu_73_in_1, msg_to_check_it_5_cnu_73_in_2, msg_to_check_it_5_cnu_73_in_3, msg_to_check_it_5_cnu_73_in_4, msg_to_check_it_5_cnu_73_in_5, msg_to_check_it_5_cnu_74_in_0, msg_to_check_it_5_cnu_74_in_1, msg_to_check_it_5_cnu_74_in_2, msg_to_check_it_5_cnu_74_in_3, msg_to_check_it_5_cnu_74_in_4, msg_to_check_it_5_cnu_74_in_5, msg_to_check_it_5_cnu_75_in_0, msg_to_check_it_5_cnu_75_in_1, msg_to_check_it_5_cnu_75_in_2, msg_to_check_it_5_cnu_75_in_3, msg_to_check_it_5_cnu_75_in_4, msg_to_check_it_5_cnu_75_in_5, msg_to_check_it_5_cnu_76_in_0, msg_to_check_it_5_cnu_76_in_1, msg_to_check_it_5_cnu_76_in_2, msg_to_check_it_5_cnu_76_in_3, msg_to_check_it_5_cnu_76_in_4, msg_to_check_it_5_cnu_76_in_5, msg_to_check_it_5_cnu_77_in_0, msg_to_check_it_5_cnu_77_in_1, msg_to_check_it_5_cnu_77_in_2, msg_to_check_it_5_cnu_77_in_3, msg_to_check_it_5_cnu_77_in_4, msg_to_check_it_5_cnu_77_in_5, msg_to_check_it_5_cnu_78_in_0, msg_to_check_it_5_cnu_78_in_1, msg_to_check_it_5_cnu_78_in_2, msg_to_check_it_5_cnu_78_in_3, msg_to_check_it_5_cnu_78_in_4, msg_to_check_it_5_cnu_78_in_5, msg_to_check_it_5_cnu_79_in_0, msg_to_check_it_5_cnu_79_in_1, msg_to_check_it_5_cnu_79_in_2, msg_to_check_it_5_cnu_79_in_3, msg_to_check_it_5_cnu_79_in_4, msg_to_check_it_5_cnu_79_in_5, msg_to_check_it_5_cnu_80_in_0, msg_to_check_it_5_cnu_80_in_1, msg_to_check_it_5_cnu_80_in_2, msg_to_check_it_5_cnu_80_in_3, msg_to_check_it_5_cnu_80_in_4, msg_to_check_it_5_cnu_80_in_5, msg_to_check_it_5_cnu_81_in_0, msg_to_check_it_5_cnu_81_in_1, msg_to_check_it_5_cnu_81_in_2, msg_to_check_it_5_cnu_81_in_3, msg_to_check_it_5_cnu_81_in_4, msg_to_check_it_5_cnu_81_in_5, msg_to_check_it_5_cnu_82_in_0, msg_to_check_it_5_cnu_82_in_1, msg_to_check_it_5_cnu_82_in_2, msg_to_check_it_5_cnu_82_in_3, msg_to_check_it_5_cnu_82_in_4, msg_to_check_it_5_cnu_82_in_5, msg_to_check_it_5_cnu_83_in_0, msg_to_check_it_5_cnu_83_in_1, msg_to_check_it_5_cnu_83_in_2, msg_to_check_it_5_cnu_83_in_3, msg_to_check_it_5_cnu_83_in_4, msg_to_check_it_5_cnu_83_in_5, msg_to_check_it_5_cnu_84_in_0, msg_to_check_it_5_cnu_84_in_1, msg_to_check_it_5_cnu_84_in_2, msg_to_check_it_5_cnu_84_in_3, msg_to_check_it_5_cnu_84_in_4, msg_to_check_it_5_cnu_84_in_5, msg_to_check_it_5_cnu_85_in_0, msg_to_check_it_5_cnu_85_in_1, msg_to_check_it_5_cnu_85_in_2, msg_to_check_it_5_cnu_85_in_3, msg_to_check_it_5_cnu_85_in_4, msg_to_check_it_5_cnu_85_in_5, msg_to_check_it_5_cnu_86_in_0, msg_to_check_it_5_cnu_86_in_1, msg_to_check_it_5_cnu_86_in_2, msg_to_check_it_5_cnu_86_in_3, msg_to_check_it_5_cnu_86_in_4, msg_to_check_it_5_cnu_86_in_5, msg_to_check_it_5_cnu_87_in_0, msg_to_check_it_5_cnu_87_in_1, msg_to_check_it_5_cnu_87_in_2, msg_to_check_it_5_cnu_87_in_3, msg_to_check_it_5_cnu_87_in_4, msg_to_check_it_5_cnu_87_in_5, msg_to_check_it_5_cnu_88_in_0, msg_to_check_it_5_cnu_88_in_1, msg_to_check_it_5_cnu_88_in_2, msg_to_check_it_5_cnu_88_in_3, msg_to_check_it_5_cnu_88_in_4, msg_to_check_it_5_cnu_88_in_5, msg_to_check_it_5_cnu_89_in_0, msg_to_check_it_5_cnu_89_in_1, msg_to_check_it_5_cnu_89_in_2, msg_to_check_it_5_cnu_89_in_3, msg_to_check_it_5_cnu_89_in_4, msg_to_check_it_5_cnu_89_in_5, msg_to_check_it_5_cnu_90_in_0, msg_to_check_it_5_cnu_90_in_1, msg_to_check_it_5_cnu_90_in_2, msg_to_check_it_5_cnu_90_in_3, msg_to_check_it_5_cnu_90_in_4, msg_to_check_it_5_cnu_90_in_5, msg_to_check_it_5_cnu_91_in_0, msg_to_check_it_5_cnu_91_in_1, msg_to_check_it_5_cnu_91_in_2, msg_to_check_it_5_cnu_91_in_3, msg_to_check_it_5_cnu_91_in_4, msg_to_check_it_5_cnu_91_in_5, msg_to_check_it_5_cnu_92_in_0, msg_to_check_it_5_cnu_92_in_1, msg_to_check_it_5_cnu_92_in_2, msg_to_check_it_5_cnu_92_in_3, msg_to_check_it_5_cnu_92_in_4, msg_to_check_it_5_cnu_92_in_5, msg_to_check_it_5_cnu_93_in_0, msg_to_check_it_5_cnu_93_in_1, msg_to_check_it_5_cnu_93_in_2, msg_to_check_it_5_cnu_93_in_3, msg_to_check_it_5_cnu_93_in_4, msg_to_check_it_5_cnu_93_in_5, msg_to_check_it_5_cnu_94_in_0, msg_to_check_it_5_cnu_94_in_1, msg_to_check_it_5_cnu_94_in_2, msg_to_check_it_5_cnu_94_in_3, msg_to_check_it_5_cnu_94_in_4, msg_to_check_it_5_cnu_94_in_5, msg_to_check_it_5_cnu_95_in_0, msg_to_check_it_5_cnu_95_in_1, msg_to_check_it_5_cnu_95_in_2, msg_to_check_it_5_cnu_95_in_3, msg_to_check_it_5_cnu_95_in_4, msg_to_check_it_5_cnu_95_in_5, msg_to_check_it_5_cnu_96_in_0, msg_to_check_it_5_cnu_96_in_1, msg_to_check_it_5_cnu_96_in_2, msg_to_check_it_5_cnu_96_in_3, msg_to_check_it_5_cnu_96_in_4, msg_to_check_it_5_cnu_96_in_5, msg_to_check_it_5_cnu_97_in_0, msg_to_check_it_5_cnu_97_in_1, msg_to_check_it_5_cnu_97_in_2, msg_to_check_it_5_cnu_97_in_3, msg_to_check_it_5_cnu_97_in_4, msg_to_check_it_5_cnu_97_in_5, msg_to_check_it_5_cnu_98_in_0, msg_to_check_it_5_cnu_98_in_1, msg_to_check_it_5_cnu_98_in_2, msg_to_check_it_5_cnu_98_in_3, msg_to_check_it_5_cnu_98_in_4, msg_to_check_it_5_cnu_98_in_5, msg_to_check_it_6_cnu_0_in_0, msg_to_check_it_6_cnu_0_in_1, msg_to_check_it_6_cnu_0_in_2, msg_to_check_it_6_cnu_0_in_3, msg_to_check_it_6_cnu_0_in_4, msg_to_check_it_6_cnu_0_in_5, msg_to_check_it_6_cnu_1_in_0, msg_to_check_it_6_cnu_1_in_1, msg_to_check_it_6_cnu_1_in_2, msg_to_check_it_6_cnu_1_in_3, msg_to_check_it_6_cnu_1_in_4, msg_to_check_it_6_cnu_1_in_5, msg_to_check_it_6_cnu_2_in_0, msg_to_check_it_6_cnu_2_in_1, msg_to_check_it_6_cnu_2_in_2, msg_to_check_it_6_cnu_2_in_3, msg_to_check_it_6_cnu_2_in_4, msg_to_check_it_6_cnu_2_in_5, msg_to_check_it_6_cnu_3_in_0, msg_to_check_it_6_cnu_3_in_1, msg_to_check_it_6_cnu_3_in_2, msg_to_check_it_6_cnu_3_in_3, msg_to_check_it_6_cnu_3_in_4, msg_to_check_it_6_cnu_3_in_5, msg_to_check_it_6_cnu_4_in_0, msg_to_check_it_6_cnu_4_in_1, msg_to_check_it_6_cnu_4_in_2, msg_to_check_it_6_cnu_4_in_3, msg_to_check_it_6_cnu_4_in_4, msg_to_check_it_6_cnu_4_in_5, msg_to_check_it_6_cnu_5_in_0, msg_to_check_it_6_cnu_5_in_1, msg_to_check_it_6_cnu_5_in_2, msg_to_check_it_6_cnu_5_in_3, msg_to_check_it_6_cnu_5_in_4, msg_to_check_it_6_cnu_5_in_5, msg_to_check_it_6_cnu_6_in_0, msg_to_check_it_6_cnu_6_in_1, msg_to_check_it_6_cnu_6_in_2, msg_to_check_it_6_cnu_6_in_3, msg_to_check_it_6_cnu_6_in_4, msg_to_check_it_6_cnu_6_in_5, msg_to_check_it_6_cnu_7_in_0, msg_to_check_it_6_cnu_7_in_1, msg_to_check_it_6_cnu_7_in_2, msg_to_check_it_6_cnu_7_in_3, msg_to_check_it_6_cnu_7_in_4, msg_to_check_it_6_cnu_7_in_5, msg_to_check_it_6_cnu_8_in_0, msg_to_check_it_6_cnu_8_in_1, msg_to_check_it_6_cnu_8_in_2, msg_to_check_it_6_cnu_8_in_3, msg_to_check_it_6_cnu_8_in_4, msg_to_check_it_6_cnu_8_in_5, msg_to_check_it_6_cnu_9_in_0, msg_to_check_it_6_cnu_9_in_1, msg_to_check_it_6_cnu_9_in_2, msg_to_check_it_6_cnu_9_in_3, msg_to_check_it_6_cnu_9_in_4, msg_to_check_it_6_cnu_9_in_5, msg_to_check_it_6_cnu_10_in_0, msg_to_check_it_6_cnu_10_in_1, msg_to_check_it_6_cnu_10_in_2, msg_to_check_it_6_cnu_10_in_3, msg_to_check_it_6_cnu_10_in_4, msg_to_check_it_6_cnu_10_in_5, msg_to_check_it_6_cnu_11_in_0, msg_to_check_it_6_cnu_11_in_1, msg_to_check_it_6_cnu_11_in_2, msg_to_check_it_6_cnu_11_in_3, msg_to_check_it_6_cnu_11_in_4, msg_to_check_it_6_cnu_11_in_5, msg_to_check_it_6_cnu_12_in_0, msg_to_check_it_6_cnu_12_in_1, msg_to_check_it_6_cnu_12_in_2, msg_to_check_it_6_cnu_12_in_3, msg_to_check_it_6_cnu_12_in_4, msg_to_check_it_6_cnu_12_in_5, msg_to_check_it_6_cnu_13_in_0, msg_to_check_it_6_cnu_13_in_1, msg_to_check_it_6_cnu_13_in_2, msg_to_check_it_6_cnu_13_in_3, msg_to_check_it_6_cnu_13_in_4, msg_to_check_it_6_cnu_13_in_5, msg_to_check_it_6_cnu_14_in_0, msg_to_check_it_6_cnu_14_in_1, msg_to_check_it_6_cnu_14_in_2, msg_to_check_it_6_cnu_14_in_3, msg_to_check_it_6_cnu_14_in_4, msg_to_check_it_6_cnu_14_in_5, msg_to_check_it_6_cnu_15_in_0, msg_to_check_it_6_cnu_15_in_1, msg_to_check_it_6_cnu_15_in_2, msg_to_check_it_6_cnu_15_in_3, msg_to_check_it_6_cnu_15_in_4, msg_to_check_it_6_cnu_15_in_5, msg_to_check_it_6_cnu_16_in_0, msg_to_check_it_6_cnu_16_in_1, msg_to_check_it_6_cnu_16_in_2, msg_to_check_it_6_cnu_16_in_3, msg_to_check_it_6_cnu_16_in_4, msg_to_check_it_6_cnu_16_in_5, msg_to_check_it_6_cnu_17_in_0, msg_to_check_it_6_cnu_17_in_1, msg_to_check_it_6_cnu_17_in_2, msg_to_check_it_6_cnu_17_in_3, msg_to_check_it_6_cnu_17_in_4, msg_to_check_it_6_cnu_17_in_5, msg_to_check_it_6_cnu_18_in_0, msg_to_check_it_6_cnu_18_in_1, msg_to_check_it_6_cnu_18_in_2, msg_to_check_it_6_cnu_18_in_3, msg_to_check_it_6_cnu_18_in_4, msg_to_check_it_6_cnu_18_in_5, msg_to_check_it_6_cnu_19_in_0, msg_to_check_it_6_cnu_19_in_1, msg_to_check_it_6_cnu_19_in_2, msg_to_check_it_6_cnu_19_in_3, msg_to_check_it_6_cnu_19_in_4, msg_to_check_it_6_cnu_19_in_5, msg_to_check_it_6_cnu_20_in_0, msg_to_check_it_6_cnu_20_in_1, msg_to_check_it_6_cnu_20_in_2, msg_to_check_it_6_cnu_20_in_3, msg_to_check_it_6_cnu_20_in_4, msg_to_check_it_6_cnu_20_in_5, msg_to_check_it_6_cnu_21_in_0, msg_to_check_it_6_cnu_21_in_1, msg_to_check_it_6_cnu_21_in_2, msg_to_check_it_6_cnu_21_in_3, msg_to_check_it_6_cnu_21_in_4, msg_to_check_it_6_cnu_21_in_5, msg_to_check_it_6_cnu_22_in_0, msg_to_check_it_6_cnu_22_in_1, msg_to_check_it_6_cnu_22_in_2, msg_to_check_it_6_cnu_22_in_3, msg_to_check_it_6_cnu_22_in_4, msg_to_check_it_6_cnu_22_in_5, msg_to_check_it_6_cnu_23_in_0, msg_to_check_it_6_cnu_23_in_1, msg_to_check_it_6_cnu_23_in_2, msg_to_check_it_6_cnu_23_in_3, msg_to_check_it_6_cnu_23_in_4, msg_to_check_it_6_cnu_23_in_5, msg_to_check_it_6_cnu_24_in_0, msg_to_check_it_6_cnu_24_in_1, msg_to_check_it_6_cnu_24_in_2, msg_to_check_it_6_cnu_24_in_3, msg_to_check_it_6_cnu_24_in_4, msg_to_check_it_6_cnu_24_in_5, msg_to_check_it_6_cnu_25_in_0, msg_to_check_it_6_cnu_25_in_1, msg_to_check_it_6_cnu_25_in_2, msg_to_check_it_6_cnu_25_in_3, msg_to_check_it_6_cnu_25_in_4, msg_to_check_it_6_cnu_25_in_5, msg_to_check_it_6_cnu_26_in_0, msg_to_check_it_6_cnu_26_in_1, msg_to_check_it_6_cnu_26_in_2, msg_to_check_it_6_cnu_26_in_3, msg_to_check_it_6_cnu_26_in_4, msg_to_check_it_6_cnu_26_in_5, msg_to_check_it_6_cnu_27_in_0, msg_to_check_it_6_cnu_27_in_1, msg_to_check_it_6_cnu_27_in_2, msg_to_check_it_6_cnu_27_in_3, msg_to_check_it_6_cnu_27_in_4, msg_to_check_it_6_cnu_27_in_5, msg_to_check_it_6_cnu_28_in_0, msg_to_check_it_6_cnu_28_in_1, msg_to_check_it_6_cnu_28_in_2, msg_to_check_it_6_cnu_28_in_3, msg_to_check_it_6_cnu_28_in_4, msg_to_check_it_6_cnu_28_in_5, msg_to_check_it_6_cnu_29_in_0, msg_to_check_it_6_cnu_29_in_1, msg_to_check_it_6_cnu_29_in_2, msg_to_check_it_6_cnu_29_in_3, msg_to_check_it_6_cnu_29_in_4, msg_to_check_it_6_cnu_29_in_5, msg_to_check_it_6_cnu_30_in_0, msg_to_check_it_6_cnu_30_in_1, msg_to_check_it_6_cnu_30_in_2, msg_to_check_it_6_cnu_30_in_3, msg_to_check_it_6_cnu_30_in_4, msg_to_check_it_6_cnu_30_in_5, msg_to_check_it_6_cnu_31_in_0, msg_to_check_it_6_cnu_31_in_1, msg_to_check_it_6_cnu_31_in_2, msg_to_check_it_6_cnu_31_in_3, msg_to_check_it_6_cnu_31_in_4, msg_to_check_it_6_cnu_31_in_5, msg_to_check_it_6_cnu_32_in_0, msg_to_check_it_6_cnu_32_in_1, msg_to_check_it_6_cnu_32_in_2, msg_to_check_it_6_cnu_32_in_3, msg_to_check_it_6_cnu_32_in_4, msg_to_check_it_6_cnu_32_in_5, msg_to_check_it_6_cnu_33_in_0, msg_to_check_it_6_cnu_33_in_1, msg_to_check_it_6_cnu_33_in_2, msg_to_check_it_6_cnu_33_in_3, msg_to_check_it_6_cnu_33_in_4, msg_to_check_it_6_cnu_33_in_5, msg_to_check_it_6_cnu_34_in_0, msg_to_check_it_6_cnu_34_in_1, msg_to_check_it_6_cnu_34_in_2, msg_to_check_it_6_cnu_34_in_3, msg_to_check_it_6_cnu_34_in_4, msg_to_check_it_6_cnu_34_in_5, msg_to_check_it_6_cnu_35_in_0, msg_to_check_it_6_cnu_35_in_1, msg_to_check_it_6_cnu_35_in_2, msg_to_check_it_6_cnu_35_in_3, msg_to_check_it_6_cnu_35_in_4, msg_to_check_it_6_cnu_35_in_5, msg_to_check_it_6_cnu_36_in_0, msg_to_check_it_6_cnu_36_in_1, msg_to_check_it_6_cnu_36_in_2, msg_to_check_it_6_cnu_36_in_3, msg_to_check_it_6_cnu_36_in_4, msg_to_check_it_6_cnu_36_in_5, msg_to_check_it_6_cnu_37_in_0, msg_to_check_it_6_cnu_37_in_1, msg_to_check_it_6_cnu_37_in_2, msg_to_check_it_6_cnu_37_in_3, msg_to_check_it_6_cnu_37_in_4, msg_to_check_it_6_cnu_37_in_5, msg_to_check_it_6_cnu_38_in_0, msg_to_check_it_6_cnu_38_in_1, msg_to_check_it_6_cnu_38_in_2, msg_to_check_it_6_cnu_38_in_3, msg_to_check_it_6_cnu_38_in_4, msg_to_check_it_6_cnu_38_in_5, msg_to_check_it_6_cnu_39_in_0, msg_to_check_it_6_cnu_39_in_1, msg_to_check_it_6_cnu_39_in_2, msg_to_check_it_6_cnu_39_in_3, msg_to_check_it_6_cnu_39_in_4, msg_to_check_it_6_cnu_39_in_5, msg_to_check_it_6_cnu_40_in_0, msg_to_check_it_6_cnu_40_in_1, msg_to_check_it_6_cnu_40_in_2, msg_to_check_it_6_cnu_40_in_3, msg_to_check_it_6_cnu_40_in_4, msg_to_check_it_6_cnu_40_in_5, msg_to_check_it_6_cnu_41_in_0, msg_to_check_it_6_cnu_41_in_1, msg_to_check_it_6_cnu_41_in_2, msg_to_check_it_6_cnu_41_in_3, msg_to_check_it_6_cnu_41_in_4, msg_to_check_it_6_cnu_41_in_5, msg_to_check_it_6_cnu_42_in_0, msg_to_check_it_6_cnu_42_in_1, msg_to_check_it_6_cnu_42_in_2, msg_to_check_it_6_cnu_42_in_3, msg_to_check_it_6_cnu_42_in_4, msg_to_check_it_6_cnu_42_in_5, msg_to_check_it_6_cnu_43_in_0, msg_to_check_it_6_cnu_43_in_1, msg_to_check_it_6_cnu_43_in_2, msg_to_check_it_6_cnu_43_in_3, msg_to_check_it_6_cnu_43_in_4, msg_to_check_it_6_cnu_43_in_5, msg_to_check_it_6_cnu_44_in_0, msg_to_check_it_6_cnu_44_in_1, msg_to_check_it_6_cnu_44_in_2, msg_to_check_it_6_cnu_44_in_3, msg_to_check_it_6_cnu_44_in_4, msg_to_check_it_6_cnu_44_in_5, msg_to_check_it_6_cnu_45_in_0, msg_to_check_it_6_cnu_45_in_1, msg_to_check_it_6_cnu_45_in_2, msg_to_check_it_6_cnu_45_in_3, msg_to_check_it_6_cnu_45_in_4, msg_to_check_it_6_cnu_45_in_5, msg_to_check_it_6_cnu_46_in_0, msg_to_check_it_6_cnu_46_in_1, msg_to_check_it_6_cnu_46_in_2, msg_to_check_it_6_cnu_46_in_3, msg_to_check_it_6_cnu_46_in_4, msg_to_check_it_6_cnu_46_in_5, msg_to_check_it_6_cnu_47_in_0, msg_to_check_it_6_cnu_47_in_1, msg_to_check_it_6_cnu_47_in_2, msg_to_check_it_6_cnu_47_in_3, msg_to_check_it_6_cnu_47_in_4, msg_to_check_it_6_cnu_47_in_5, msg_to_check_it_6_cnu_48_in_0, msg_to_check_it_6_cnu_48_in_1, msg_to_check_it_6_cnu_48_in_2, msg_to_check_it_6_cnu_48_in_3, msg_to_check_it_6_cnu_48_in_4, msg_to_check_it_6_cnu_48_in_5, msg_to_check_it_6_cnu_49_in_0, msg_to_check_it_6_cnu_49_in_1, msg_to_check_it_6_cnu_49_in_2, msg_to_check_it_6_cnu_49_in_3, msg_to_check_it_6_cnu_49_in_4, msg_to_check_it_6_cnu_49_in_5, msg_to_check_it_6_cnu_50_in_0, msg_to_check_it_6_cnu_50_in_1, msg_to_check_it_6_cnu_50_in_2, msg_to_check_it_6_cnu_50_in_3, msg_to_check_it_6_cnu_50_in_4, msg_to_check_it_6_cnu_50_in_5, msg_to_check_it_6_cnu_51_in_0, msg_to_check_it_6_cnu_51_in_1, msg_to_check_it_6_cnu_51_in_2, msg_to_check_it_6_cnu_51_in_3, msg_to_check_it_6_cnu_51_in_4, msg_to_check_it_6_cnu_51_in_5, msg_to_check_it_6_cnu_52_in_0, msg_to_check_it_6_cnu_52_in_1, msg_to_check_it_6_cnu_52_in_2, msg_to_check_it_6_cnu_52_in_3, msg_to_check_it_6_cnu_52_in_4, msg_to_check_it_6_cnu_52_in_5, msg_to_check_it_6_cnu_53_in_0, msg_to_check_it_6_cnu_53_in_1, msg_to_check_it_6_cnu_53_in_2, msg_to_check_it_6_cnu_53_in_3, msg_to_check_it_6_cnu_53_in_4, msg_to_check_it_6_cnu_53_in_5, msg_to_check_it_6_cnu_54_in_0, msg_to_check_it_6_cnu_54_in_1, msg_to_check_it_6_cnu_54_in_2, msg_to_check_it_6_cnu_54_in_3, msg_to_check_it_6_cnu_54_in_4, msg_to_check_it_6_cnu_54_in_5, msg_to_check_it_6_cnu_55_in_0, msg_to_check_it_6_cnu_55_in_1, msg_to_check_it_6_cnu_55_in_2, msg_to_check_it_6_cnu_55_in_3, msg_to_check_it_6_cnu_55_in_4, msg_to_check_it_6_cnu_55_in_5, msg_to_check_it_6_cnu_56_in_0, msg_to_check_it_6_cnu_56_in_1, msg_to_check_it_6_cnu_56_in_2, msg_to_check_it_6_cnu_56_in_3, msg_to_check_it_6_cnu_56_in_4, msg_to_check_it_6_cnu_56_in_5, msg_to_check_it_6_cnu_57_in_0, msg_to_check_it_6_cnu_57_in_1, msg_to_check_it_6_cnu_57_in_2, msg_to_check_it_6_cnu_57_in_3, msg_to_check_it_6_cnu_57_in_4, msg_to_check_it_6_cnu_57_in_5, msg_to_check_it_6_cnu_58_in_0, msg_to_check_it_6_cnu_58_in_1, msg_to_check_it_6_cnu_58_in_2, msg_to_check_it_6_cnu_58_in_3, msg_to_check_it_6_cnu_58_in_4, msg_to_check_it_6_cnu_58_in_5, msg_to_check_it_6_cnu_59_in_0, msg_to_check_it_6_cnu_59_in_1, msg_to_check_it_6_cnu_59_in_2, msg_to_check_it_6_cnu_59_in_3, msg_to_check_it_6_cnu_59_in_4, msg_to_check_it_6_cnu_59_in_5, msg_to_check_it_6_cnu_60_in_0, msg_to_check_it_6_cnu_60_in_1, msg_to_check_it_6_cnu_60_in_2, msg_to_check_it_6_cnu_60_in_3, msg_to_check_it_6_cnu_60_in_4, msg_to_check_it_6_cnu_60_in_5, msg_to_check_it_6_cnu_61_in_0, msg_to_check_it_6_cnu_61_in_1, msg_to_check_it_6_cnu_61_in_2, msg_to_check_it_6_cnu_61_in_3, msg_to_check_it_6_cnu_61_in_4, msg_to_check_it_6_cnu_61_in_5, msg_to_check_it_6_cnu_62_in_0, msg_to_check_it_6_cnu_62_in_1, msg_to_check_it_6_cnu_62_in_2, msg_to_check_it_6_cnu_62_in_3, msg_to_check_it_6_cnu_62_in_4, msg_to_check_it_6_cnu_62_in_5, msg_to_check_it_6_cnu_63_in_0, msg_to_check_it_6_cnu_63_in_1, msg_to_check_it_6_cnu_63_in_2, msg_to_check_it_6_cnu_63_in_3, msg_to_check_it_6_cnu_63_in_4, msg_to_check_it_6_cnu_63_in_5, msg_to_check_it_6_cnu_64_in_0, msg_to_check_it_6_cnu_64_in_1, msg_to_check_it_6_cnu_64_in_2, msg_to_check_it_6_cnu_64_in_3, msg_to_check_it_6_cnu_64_in_4, msg_to_check_it_6_cnu_64_in_5, msg_to_check_it_6_cnu_65_in_0, msg_to_check_it_6_cnu_65_in_1, msg_to_check_it_6_cnu_65_in_2, msg_to_check_it_6_cnu_65_in_3, msg_to_check_it_6_cnu_65_in_4, msg_to_check_it_6_cnu_65_in_5, msg_to_check_it_6_cnu_66_in_0, msg_to_check_it_6_cnu_66_in_1, msg_to_check_it_6_cnu_66_in_2, msg_to_check_it_6_cnu_66_in_3, msg_to_check_it_6_cnu_66_in_4, msg_to_check_it_6_cnu_66_in_5, msg_to_check_it_6_cnu_67_in_0, msg_to_check_it_6_cnu_67_in_1, msg_to_check_it_6_cnu_67_in_2, msg_to_check_it_6_cnu_67_in_3, msg_to_check_it_6_cnu_67_in_4, msg_to_check_it_6_cnu_67_in_5, msg_to_check_it_6_cnu_68_in_0, msg_to_check_it_6_cnu_68_in_1, msg_to_check_it_6_cnu_68_in_2, msg_to_check_it_6_cnu_68_in_3, msg_to_check_it_6_cnu_68_in_4, msg_to_check_it_6_cnu_68_in_5, msg_to_check_it_6_cnu_69_in_0, msg_to_check_it_6_cnu_69_in_1, msg_to_check_it_6_cnu_69_in_2, msg_to_check_it_6_cnu_69_in_3, msg_to_check_it_6_cnu_69_in_4, msg_to_check_it_6_cnu_69_in_5, msg_to_check_it_6_cnu_70_in_0, msg_to_check_it_6_cnu_70_in_1, msg_to_check_it_6_cnu_70_in_2, msg_to_check_it_6_cnu_70_in_3, msg_to_check_it_6_cnu_70_in_4, msg_to_check_it_6_cnu_70_in_5, msg_to_check_it_6_cnu_71_in_0, msg_to_check_it_6_cnu_71_in_1, msg_to_check_it_6_cnu_71_in_2, msg_to_check_it_6_cnu_71_in_3, msg_to_check_it_6_cnu_71_in_4, msg_to_check_it_6_cnu_71_in_5, msg_to_check_it_6_cnu_72_in_0, msg_to_check_it_6_cnu_72_in_1, msg_to_check_it_6_cnu_72_in_2, msg_to_check_it_6_cnu_72_in_3, msg_to_check_it_6_cnu_72_in_4, msg_to_check_it_6_cnu_72_in_5, msg_to_check_it_6_cnu_73_in_0, msg_to_check_it_6_cnu_73_in_1, msg_to_check_it_6_cnu_73_in_2, msg_to_check_it_6_cnu_73_in_3, msg_to_check_it_6_cnu_73_in_4, msg_to_check_it_6_cnu_73_in_5, msg_to_check_it_6_cnu_74_in_0, msg_to_check_it_6_cnu_74_in_1, msg_to_check_it_6_cnu_74_in_2, msg_to_check_it_6_cnu_74_in_3, msg_to_check_it_6_cnu_74_in_4, msg_to_check_it_6_cnu_74_in_5, msg_to_check_it_6_cnu_75_in_0, msg_to_check_it_6_cnu_75_in_1, msg_to_check_it_6_cnu_75_in_2, msg_to_check_it_6_cnu_75_in_3, msg_to_check_it_6_cnu_75_in_4, msg_to_check_it_6_cnu_75_in_5, msg_to_check_it_6_cnu_76_in_0, msg_to_check_it_6_cnu_76_in_1, msg_to_check_it_6_cnu_76_in_2, msg_to_check_it_6_cnu_76_in_3, msg_to_check_it_6_cnu_76_in_4, msg_to_check_it_6_cnu_76_in_5, msg_to_check_it_6_cnu_77_in_0, msg_to_check_it_6_cnu_77_in_1, msg_to_check_it_6_cnu_77_in_2, msg_to_check_it_6_cnu_77_in_3, msg_to_check_it_6_cnu_77_in_4, msg_to_check_it_6_cnu_77_in_5, msg_to_check_it_6_cnu_78_in_0, msg_to_check_it_6_cnu_78_in_1, msg_to_check_it_6_cnu_78_in_2, msg_to_check_it_6_cnu_78_in_3, msg_to_check_it_6_cnu_78_in_4, msg_to_check_it_6_cnu_78_in_5, msg_to_check_it_6_cnu_79_in_0, msg_to_check_it_6_cnu_79_in_1, msg_to_check_it_6_cnu_79_in_2, msg_to_check_it_6_cnu_79_in_3, msg_to_check_it_6_cnu_79_in_4, msg_to_check_it_6_cnu_79_in_5, msg_to_check_it_6_cnu_80_in_0, msg_to_check_it_6_cnu_80_in_1, msg_to_check_it_6_cnu_80_in_2, msg_to_check_it_6_cnu_80_in_3, msg_to_check_it_6_cnu_80_in_4, msg_to_check_it_6_cnu_80_in_5, msg_to_check_it_6_cnu_81_in_0, msg_to_check_it_6_cnu_81_in_1, msg_to_check_it_6_cnu_81_in_2, msg_to_check_it_6_cnu_81_in_3, msg_to_check_it_6_cnu_81_in_4, msg_to_check_it_6_cnu_81_in_5, msg_to_check_it_6_cnu_82_in_0, msg_to_check_it_6_cnu_82_in_1, msg_to_check_it_6_cnu_82_in_2, msg_to_check_it_6_cnu_82_in_3, msg_to_check_it_6_cnu_82_in_4, msg_to_check_it_6_cnu_82_in_5, msg_to_check_it_6_cnu_83_in_0, msg_to_check_it_6_cnu_83_in_1, msg_to_check_it_6_cnu_83_in_2, msg_to_check_it_6_cnu_83_in_3, msg_to_check_it_6_cnu_83_in_4, msg_to_check_it_6_cnu_83_in_5, msg_to_check_it_6_cnu_84_in_0, msg_to_check_it_6_cnu_84_in_1, msg_to_check_it_6_cnu_84_in_2, msg_to_check_it_6_cnu_84_in_3, msg_to_check_it_6_cnu_84_in_4, msg_to_check_it_6_cnu_84_in_5, msg_to_check_it_6_cnu_85_in_0, msg_to_check_it_6_cnu_85_in_1, msg_to_check_it_6_cnu_85_in_2, msg_to_check_it_6_cnu_85_in_3, msg_to_check_it_6_cnu_85_in_4, msg_to_check_it_6_cnu_85_in_5, msg_to_check_it_6_cnu_86_in_0, msg_to_check_it_6_cnu_86_in_1, msg_to_check_it_6_cnu_86_in_2, msg_to_check_it_6_cnu_86_in_3, msg_to_check_it_6_cnu_86_in_4, msg_to_check_it_6_cnu_86_in_5, msg_to_check_it_6_cnu_87_in_0, msg_to_check_it_6_cnu_87_in_1, msg_to_check_it_6_cnu_87_in_2, msg_to_check_it_6_cnu_87_in_3, msg_to_check_it_6_cnu_87_in_4, msg_to_check_it_6_cnu_87_in_5, msg_to_check_it_6_cnu_88_in_0, msg_to_check_it_6_cnu_88_in_1, msg_to_check_it_6_cnu_88_in_2, msg_to_check_it_6_cnu_88_in_3, msg_to_check_it_6_cnu_88_in_4, msg_to_check_it_6_cnu_88_in_5, msg_to_check_it_6_cnu_89_in_0, msg_to_check_it_6_cnu_89_in_1, msg_to_check_it_6_cnu_89_in_2, msg_to_check_it_6_cnu_89_in_3, msg_to_check_it_6_cnu_89_in_4, msg_to_check_it_6_cnu_89_in_5, msg_to_check_it_6_cnu_90_in_0, msg_to_check_it_6_cnu_90_in_1, msg_to_check_it_6_cnu_90_in_2, msg_to_check_it_6_cnu_90_in_3, msg_to_check_it_6_cnu_90_in_4, msg_to_check_it_6_cnu_90_in_5, msg_to_check_it_6_cnu_91_in_0, msg_to_check_it_6_cnu_91_in_1, msg_to_check_it_6_cnu_91_in_2, msg_to_check_it_6_cnu_91_in_3, msg_to_check_it_6_cnu_91_in_4, msg_to_check_it_6_cnu_91_in_5, msg_to_check_it_6_cnu_92_in_0, msg_to_check_it_6_cnu_92_in_1, msg_to_check_it_6_cnu_92_in_2, msg_to_check_it_6_cnu_92_in_3, msg_to_check_it_6_cnu_92_in_4, msg_to_check_it_6_cnu_92_in_5, msg_to_check_it_6_cnu_93_in_0, msg_to_check_it_6_cnu_93_in_1, msg_to_check_it_6_cnu_93_in_2, msg_to_check_it_6_cnu_93_in_3, msg_to_check_it_6_cnu_93_in_4, msg_to_check_it_6_cnu_93_in_5, msg_to_check_it_6_cnu_94_in_0, msg_to_check_it_6_cnu_94_in_1, msg_to_check_it_6_cnu_94_in_2, msg_to_check_it_6_cnu_94_in_3, msg_to_check_it_6_cnu_94_in_4, msg_to_check_it_6_cnu_94_in_5, msg_to_check_it_6_cnu_95_in_0, msg_to_check_it_6_cnu_95_in_1, msg_to_check_it_6_cnu_95_in_2, msg_to_check_it_6_cnu_95_in_3, msg_to_check_it_6_cnu_95_in_4, msg_to_check_it_6_cnu_95_in_5, msg_to_check_it_6_cnu_96_in_0, msg_to_check_it_6_cnu_96_in_1, msg_to_check_it_6_cnu_96_in_2, msg_to_check_it_6_cnu_96_in_3, msg_to_check_it_6_cnu_96_in_4, msg_to_check_it_6_cnu_96_in_5, msg_to_check_it_6_cnu_97_in_0, msg_to_check_it_6_cnu_97_in_1, msg_to_check_it_6_cnu_97_in_2, msg_to_check_it_6_cnu_97_in_3, msg_to_check_it_6_cnu_97_in_4, msg_to_check_it_6_cnu_97_in_5, msg_to_check_it_6_cnu_98_in_0, msg_to_check_it_6_cnu_98_in_1, msg_to_check_it_6_cnu_98_in_2, msg_to_check_it_6_cnu_98_in_3, msg_to_check_it_6_cnu_98_in_4, msg_to_check_it_6_cnu_98_in_5, msg_to_check_it_7_cnu_0_in_0, msg_to_check_it_7_cnu_0_in_1, msg_to_check_it_7_cnu_0_in_2, msg_to_check_it_7_cnu_0_in_3, msg_to_check_it_7_cnu_0_in_4, msg_to_check_it_7_cnu_0_in_5, msg_to_check_it_7_cnu_1_in_0, msg_to_check_it_7_cnu_1_in_1, msg_to_check_it_7_cnu_1_in_2, msg_to_check_it_7_cnu_1_in_3, msg_to_check_it_7_cnu_1_in_4, msg_to_check_it_7_cnu_1_in_5, msg_to_check_it_7_cnu_2_in_0, msg_to_check_it_7_cnu_2_in_1, msg_to_check_it_7_cnu_2_in_2, msg_to_check_it_7_cnu_2_in_3, msg_to_check_it_7_cnu_2_in_4, msg_to_check_it_7_cnu_2_in_5, msg_to_check_it_7_cnu_3_in_0, msg_to_check_it_7_cnu_3_in_1, msg_to_check_it_7_cnu_3_in_2, msg_to_check_it_7_cnu_3_in_3, msg_to_check_it_7_cnu_3_in_4, msg_to_check_it_7_cnu_3_in_5, msg_to_check_it_7_cnu_4_in_0, msg_to_check_it_7_cnu_4_in_1, msg_to_check_it_7_cnu_4_in_2, msg_to_check_it_7_cnu_4_in_3, msg_to_check_it_7_cnu_4_in_4, msg_to_check_it_7_cnu_4_in_5, msg_to_check_it_7_cnu_5_in_0, msg_to_check_it_7_cnu_5_in_1, msg_to_check_it_7_cnu_5_in_2, msg_to_check_it_7_cnu_5_in_3, msg_to_check_it_7_cnu_5_in_4, msg_to_check_it_7_cnu_5_in_5, msg_to_check_it_7_cnu_6_in_0, msg_to_check_it_7_cnu_6_in_1, msg_to_check_it_7_cnu_6_in_2, msg_to_check_it_7_cnu_6_in_3, msg_to_check_it_7_cnu_6_in_4, msg_to_check_it_7_cnu_6_in_5, msg_to_check_it_7_cnu_7_in_0, msg_to_check_it_7_cnu_7_in_1, msg_to_check_it_7_cnu_7_in_2, msg_to_check_it_7_cnu_7_in_3, msg_to_check_it_7_cnu_7_in_4, msg_to_check_it_7_cnu_7_in_5, msg_to_check_it_7_cnu_8_in_0, msg_to_check_it_7_cnu_8_in_1, msg_to_check_it_7_cnu_8_in_2, msg_to_check_it_7_cnu_8_in_3, msg_to_check_it_7_cnu_8_in_4, msg_to_check_it_7_cnu_8_in_5, msg_to_check_it_7_cnu_9_in_0, msg_to_check_it_7_cnu_9_in_1, msg_to_check_it_7_cnu_9_in_2, msg_to_check_it_7_cnu_9_in_3, msg_to_check_it_7_cnu_9_in_4, msg_to_check_it_7_cnu_9_in_5, msg_to_check_it_7_cnu_10_in_0, msg_to_check_it_7_cnu_10_in_1, msg_to_check_it_7_cnu_10_in_2, msg_to_check_it_7_cnu_10_in_3, msg_to_check_it_7_cnu_10_in_4, msg_to_check_it_7_cnu_10_in_5, msg_to_check_it_7_cnu_11_in_0, msg_to_check_it_7_cnu_11_in_1, msg_to_check_it_7_cnu_11_in_2, msg_to_check_it_7_cnu_11_in_3, msg_to_check_it_7_cnu_11_in_4, msg_to_check_it_7_cnu_11_in_5, msg_to_check_it_7_cnu_12_in_0, msg_to_check_it_7_cnu_12_in_1, msg_to_check_it_7_cnu_12_in_2, msg_to_check_it_7_cnu_12_in_3, msg_to_check_it_7_cnu_12_in_4, msg_to_check_it_7_cnu_12_in_5, msg_to_check_it_7_cnu_13_in_0, msg_to_check_it_7_cnu_13_in_1, msg_to_check_it_7_cnu_13_in_2, msg_to_check_it_7_cnu_13_in_3, msg_to_check_it_7_cnu_13_in_4, msg_to_check_it_7_cnu_13_in_5, msg_to_check_it_7_cnu_14_in_0, msg_to_check_it_7_cnu_14_in_1, msg_to_check_it_7_cnu_14_in_2, msg_to_check_it_7_cnu_14_in_3, msg_to_check_it_7_cnu_14_in_4, msg_to_check_it_7_cnu_14_in_5, msg_to_check_it_7_cnu_15_in_0, msg_to_check_it_7_cnu_15_in_1, msg_to_check_it_7_cnu_15_in_2, msg_to_check_it_7_cnu_15_in_3, msg_to_check_it_7_cnu_15_in_4, msg_to_check_it_7_cnu_15_in_5, msg_to_check_it_7_cnu_16_in_0, msg_to_check_it_7_cnu_16_in_1, msg_to_check_it_7_cnu_16_in_2, msg_to_check_it_7_cnu_16_in_3, msg_to_check_it_7_cnu_16_in_4, msg_to_check_it_7_cnu_16_in_5, msg_to_check_it_7_cnu_17_in_0, msg_to_check_it_7_cnu_17_in_1, msg_to_check_it_7_cnu_17_in_2, msg_to_check_it_7_cnu_17_in_3, msg_to_check_it_7_cnu_17_in_4, msg_to_check_it_7_cnu_17_in_5, msg_to_check_it_7_cnu_18_in_0, msg_to_check_it_7_cnu_18_in_1, msg_to_check_it_7_cnu_18_in_2, msg_to_check_it_7_cnu_18_in_3, msg_to_check_it_7_cnu_18_in_4, msg_to_check_it_7_cnu_18_in_5, msg_to_check_it_7_cnu_19_in_0, msg_to_check_it_7_cnu_19_in_1, msg_to_check_it_7_cnu_19_in_2, msg_to_check_it_7_cnu_19_in_3, msg_to_check_it_7_cnu_19_in_4, msg_to_check_it_7_cnu_19_in_5, msg_to_check_it_7_cnu_20_in_0, msg_to_check_it_7_cnu_20_in_1, msg_to_check_it_7_cnu_20_in_2, msg_to_check_it_7_cnu_20_in_3, msg_to_check_it_7_cnu_20_in_4, msg_to_check_it_7_cnu_20_in_5, msg_to_check_it_7_cnu_21_in_0, msg_to_check_it_7_cnu_21_in_1, msg_to_check_it_7_cnu_21_in_2, msg_to_check_it_7_cnu_21_in_3, msg_to_check_it_7_cnu_21_in_4, msg_to_check_it_7_cnu_21_in_5, msg_to_check_it_7_cnu_22_in_0, msg_to_check_it_7_cnu_22_in_1, msg_to_check_it_7_cnu_22_in_2, msg_to_check_it_7_cnu_22_in_3, msg_to_check_it_7_cnu_22_in_4, msg_to_check_it_7_cnu_22_in_5, msg_to_check_it_7_cnu_23_in_0, msg_to_check_it_7_cnu_23_in_1, msg_to_check_it_7_cnu_23_in_2, msg_to_check_it_7_cnu_23_in_3, msg_to_check_it_7_cnu_23_in_4, msg_to_check_it_7_cnu_23_in_5, msg_to_check_it_7_cnu_24_in_0, msg_to_check_it_7_cnu_24_in_1, msg_to_check_it_7_cnu_24_in_2, msg_to_check_it_7_cnu_24_in_3, msg_to_check_it_7_cnu_24_in_4, msg_to_check_it_7_cnu_24_in_5, msg_to_check_it_7_cnu_25_in_0, msg_to_check_it_7_cnu_25_in_1, msg_to_check_it_7_cnu_25_in_2, msg_to_check_it_7_cnu_25_in_3, msg_to_check_it_7_cnu_25_in_4, msg_to_check_it_7_cnu_25_in_5, msg_to_check_it_7_cnu_26_in_0, msg_to_check_it_7_cnu_26_in_1, msg_to_check_it_7_cnu_26_in_2, msg_to_check_it_7_cnu_26_in_3, msg_to_check_it_7_cnu_26_in_4, msg_to_check_it_7_cnu_26_in_5, msg_to_check_it_7_cnu_27_in_0, msg_to_check_it_7_cnu_27_in_1, msg_to_check_it_7_cnu_27_in_2, msg_to_check_it_7_cnu_27_in_3, msg_to_check_it_7_cnu_27_in_4, msg_to_check_it_7_cnu_27_in_5, msg_to_check_it_7_cnu_28_in_0, msg_to_check_it_7_cnu_28_in_1, msg_to_check_it_7_cnu_28_in_2, msg_to_check_it_7_cnu_28_in_3, msg_to_check_it_7_cnu_28_in_4, msg_to_check_it_7_cnu_28_in_5, msg_to_check_it_7_cnu_29_in_0, msg_to_check_it_7_cnu_29_in_1, msg_to_check_it_7_cnu_29_in_2, msg_to_check_it_7_cnu_29_in_3, msg_to_check_it_7_cnu_29_in_4, msg_to_check_it_7_cnu_29_in_5, msg_to_check_it_7_cnu_30_in_0, msg_to_check_it_7_cnu_30_in_1, msg_to_check_it_7_cnu_30_in_2, msg_to_check_it_7_cnu_30_in_3, msg_to_check_it_7_cnu_30_in_4, msg_to_check_it_7_cnu_30_in_5, msg_to_check_it_7_cnu_31_in_0, msg_to_check_it_7_cnu_31_in_1, msg_to_check_it_7_cnu_31_in_2, msg_to_check_it_7_cnu_31_in_3, msg_to_check_it_7_cnu_31_in_4, msg_to_check_it_7_cnu_31_in_5, msg_to_check_it_7_cnu_32_in_0, msg_to_check_it_7_cnu_32_in_1, msg_to_check_it_7_cnu_32_in_2, msg_to_check_it_7_cnu_32_in_3, msg_to_check_it_7_cnu_32_in_4, msg_to_check_it_7_cnu_32_in_5, msg_to_check_it_7_cnu_33_in_0, msg_to_check_it_7_cnu_33_in_1, msg_to_check_it_7_cnu_33_in_2, msg_to_check_it_7_cnu_33_in_3, msg_to_check_it_7_cnu_33_in_4, msg_to_check_it_7_cnu_33_in_5, msg_to_check_it_7_cnu_34_in_0, msg_to_check_it_7_cnu_34_in_1, msg_to_check_it_7_cnu_34_in_2, msg_to_check_it_7_cnu_34_in_3, msg_to_check_it_7_cnu_34_in_4, msg_to_check_it_7_cnu_34_in_5, msg_to_check_it_7_cnu_35_in_0, msg_to_check_it_7_cnu_35_in_1, msg_to_check_it_7_cnu_35_in_2, msg_to_check_it_7_cnu_35_in_3, msg_to_check_it_7_cnu_35_in_4, msg_to_check_it_7_cnu_35_in_5, msg_to_check_it_7_cnu_36_in_0, msg_to_check_it_7_cnu_36_in_1, msg_to_check_it_7_cnu_36_in_2, msg_to_check_it_7_cnu_36_in_3, msg_to_check_it_7_cnu_36_in_4, msg_to_check_it_7_cnu_36_in_5, msg_to_check_it_7_cnu_37_in_0, msg_to_check_it_7_cnu_37_in_1, msg_to_check_it_7_cnu_37_in_2, msg_to_check_it_7_cnu_37_in_3, msg_to_check_it_7_cnu_37_in_4, msg_to_check_it_7_cnu_37_in_5, msg_to_check_it_7_cnu_38_in_0, msg_to_check_it_7_cnu_38_in_1, msg_to_check_it_7_cnu_38_in_2, msg_to_check_it_7_cnu_38_in_3, msg_to_check_it_7_cnu_38_in_4, msg_to_check_it_7_cnu_38_in_5, msg_to_check_it_7_cnu_39_in_0, msg_to_check_it_7_cnu_39_in_1, msg_to_check_it_7_cnu_39_in_2, msg_to_check_it_7_cnu_39_in_3, msg_to_check_it_7_cnu_39_in_4, msg_to_check_it_7_cnu_39_in_5, msg_to_check_it_7_cnu_40_in_0, msg_to_check_it_7_cnu_40_in_1, msg_to_check_it_7_cnu_40_in_2, msg_to_check_it_7_cnu_40_in_3, msg_to_check_it_7_cnu_40_in_4, msg_to_check_it_7_cnu_40_in_5, msg_to_check_it_7_cnu_41_in_0, msg_to_check_it_7_cnu_41_in_1, msg_to_check_it_7_cnu_41_in_2, msg_to_check_it_7_cnu_41_in_3, msg_to_check_it_7_cnu_41_in_4, msg_to_check_it_7_cnu_41_in_5, msg_to_check_it_7_cnu_42_in_0, msg_to_check_it_7_cnu_42_in_1, msg_to_check_it_7_cnu_42_in_2, msg_to_check_it_7_cnu_42_in_3, msg_to_check_it_7_cnu_42_in_4, msg_to_check_it_7_cnu_42_in_5, msg_to_check_it_7_cnu_43_in_0, msg_to_check_it_7_cnu_43_in_1, msg_to_check_it_7_cnu_43_in_2, msg_to_check_it_7_cnu_43_in_3, msg_to_check_it_7_cnu_43_in_4, msg_to_check_it_7_cnu_43_in_5, msg_to_check_it_7_cnu_44_in_0, msg_to_check_it_7_cnu_44_in_1, msg_to_check_it_7_cnu_44_in_2, msg_to_check_it_7_cnu_44_in_3, msg_to_check_it_7_cnu_44_in_4, msg_to_check_it_7_cnu_44_in_5, msg_to_check_it_7_cnu_45_in_0, msg_to_check_it_7_cnu_45_in_1, msg_to_check_it_7_cnu_45_in_2, msg_to_check_it_7_cnu_45_in_3, msg_to_check_it_7_cnu_45_in_4, msg_to_check_it_7_cnu_45_in_5, msg_to_check_it_7_cnu_46_in_0, msg_to_check_it_7_cnu_46_in_1, msg_to_check_it_7_cnu_46_in_2, msg_to_check_it_7_cnu_46_in_3, msg_to_check_it_7_cnu_46_in_4, msg_to_check_it_7_cnu_46_in_5, msg_to_check_it_7_cnu_47_in_0, msg_to_check_it_7_cnu_47_in_1, msg_to_check_it_7_cnu_47_in_2, msg_to_check_it_7_cnu_47_in_3, msg_to_check_it_7_cnu_47_in_4, msg_to_check_it_7_cnu_47_in_5, msg_to_check_it_7_cnu_48_in_0, msg_to_check_it_7_cnu_48_in_1, msg_to_check_it_7_cnu_48_in_2, msg_to_check_it_7_cnu_48_in_3, msg_to_check_it_7_cnu_48_in_4, msg_to_check_it_7_cnu_48_in_5, msg_to_check_it_7_cnu_49_in_0, msg_to_check_it_7_cnu_49_in_1, msg_to_check_it_7_cnu_49_in_2, msg_to_check_it_7_cnu_49_in_3, msg_to_check_it_7_cnu_49_in_4, msg_to_check_it_7_cnu_49_in_5, msg_to_check_it_7_cnu_50_in_0, msg_to_check_it_7_cnu_50_in_1, msg_to_check_it_7_cnu_50_in_2, msg_to_check_it_7_cnu_50_in_3, msg_to_check_it_7_cnu_50_in_4, msg_to_check_it_7_cnu_50_in_5, msg_to_check_it_7_cnu_51_in_0, msg_to_check_it_7_cnu_51_in_1, msg_to_check_it_7_cnu_51_in_2, msg_to_check_it_7_cnu_51_in_3, msg_to_check_it_7_cnu_51_in_4, msg_to_check_it_7_cnu_51_in_5, msg_to_check_it_7_cnu_52_in_0, msg_to_check_it_7_cnu_52_in_1, msg_to_check_it_7_cnu_52_in_2, msg_to_check_it_7_cnu_52_in_3, msg_to_check_it_7_cnu_52_in_4, msg_to_check_it_7_cnu_52_in_5, msg_to_check_it_7_cnu_53_in_0, msg_to_check_it_7_cnu_53_in_1, msg_to_check_it_7_cnu_53_in_2, msg_to_check_it_7_cnu_53_in_3, msg_to_check_it_7_cnu_53_in_4, msg_to_check_it_7_cnu_53_in_5, msg_to_check_it_7_cnu_54_in_0, msg_to_check_it_7_cnu_54_in_1, msg_to_check_it_7_cnu_54_in_2, msg_to_check_it_7_cnu_54_in_3, msg_to_check_it_7_cnu_54_in_4, msg_to_check_it_7_cnu_54_in_5, msg_to_check_it_7_cnu_55_in_0, msg_to_check_it_7_cnu_55_in_1, msg_to_check_it_7_cnu_55_in_2, msg_to_check_it_7_cnu_55_in_3, msg_to_check_it_7_cnu_55_in_4, msg_to_check_it_7_cnu_55_in_5, msg_to_check_it_7_cnu_56_in_0, msg_to_check_it_7_cnu_56_in_1, msg_to_check_it_7_cnu_56_in_2, msg_to_check_it_7_cnu_56_in_3, msg_to_check_it_7_cnu_56_in_4, msg_to_check_it_7_cnu_56_in_5, msg_to_check_it_7_cnu_57_in_0, msg_to_check_it_7_cnu_57_in_1, msg_to_check_it_7_cnu_57_in_2, msg_to_check_it_7_cnu_57_in_3, msg_to_check_it_7_cnu_57_in_4, msg_to_check_it_7_cnu_57_in_5, msg_to_check_it_7_cnu_58_in_0, msg_to_check_it_7_cnu_58_in_1, msg_to_check_it_7_cnu_58_in_2, msg_to_check_it_7_cnu_58_in_3, msg_to_check_it_7_cnu_58_in_4, msg_to_check_it_7_cnu_58_in_5, msg_to_check_it_7_cnu_59_in_0, msg_to_check_it_7_cnu_59_in_1, msg_to_check_it_7_cnu_59_in_2, msg_to_check_it_7_cnu_59_in_3, msg_to_check_it_7_cnu_59_in_4, msg_to_check_it_7_cnu_59_in_5, msg_to_check_it_7_cnu_60_in_0, msg_to_check_it_7_cnu_60_in_1, msg_to_check_it_7_cnu_60_in_2, msg_to_check_it_7_cnu_60_in_3, msg_to_check_it_7_cnu_60_in_4, msg_to_check_it_7_cnu_60_in_5, msg_to_check_it_7_cnu_61_in_0, msg_to_check_it_7_cnu_61_in_1, msg_to_check_it_7_cnu_61_in_2, msg_to_check_it_7_cnu_61_in_3, msg_to_check_it_7_cnu_61_in_4, msg_to_check_it_7_cnu_61_in_5, msg_to_check_it_7_cnu_62_in_0, msg_to_check_it_7_cnu_62_in_1, msg_to_check_it_7_cnu_62_in_2, msg_to_check_it_7_cnu_62_in_3, msg_to_check_it_7_cnu_62_in_4, msg_to_check_it_7_cnu_62_in_5, msg_to_check_it_7_cnu_63_in_0, msg_to_check_it_7_cnu_63_in_1, msg_to_check_it_7_cnu_63_in_2, msg_to_check_it_7_cnu_63_in_3, msg_to_check_it_7_cnu_63_in_4, msg_to_check_it_7_cnu_63_in_5, msg_to_check_it_7_cnu_64_in_0, msg_to_check_it_7_cnu_64_in_1, msg_to_check_it_7_cnu_64_in_2, msg_to_check_it_7_cnu_64_in_3, msg_to_check_it_7_cnu_64_in_4, msg_to_check_it_7_cnu_64_in_5, msg_to_check_it_7_cnu_65_in_0, msg_to_check_it_7_cnu_65_in_1, msg_to_check_it_7_cnu_65_in_2, msg_to_check_it_7_cnu_65_in_3, msg_to_check_it_7_cnu_65_in_4, msg_to_check_it_7_cnu_65_in_5, msg_to_check_it_7_cnu_66_in_0, msg_to_check_it_7_cnu_66_in_1, msg_to_check_it_7_cnu_66_in_2, msg_to_check_it_7_cnu_66_in_3, msg_to_check_it_7_cnu_66_in_4, msg_to_check_it_7_cnu_66_in_5, msg_to_check_it_7_cnu_67_in_0, msg_to_check_it_7_cnu_67_in_1, msg_to_check_it_7_cnu_67_in_2, msg_to_check_it_7_cnu_67_in_3, msg_to_check_it_7_cnu_67_in_4, msg_to_check_it_7_cnu_67_in_5, msg_to_check_it_7_cnu_68_in_0, msg_to_check_it_7_cnu_68_in_1, msg_to_check_it_7_cnu_68_in_2, msg_to_check_it_7_cnu_68_in_3, msg_to_check_it_7_cnu_68_in_4, msg_to_check_it_7_cnu_68_in_5, msg_to_check_it_7_cnu_69_in_0, msg_to_check_it_7_cnu_69_in_1, msg_to_check_it_7_cnu_69_in_2, msg_to_check_it_7_cnu_69_in_3, msg_to_check_it_7_cnu_69_in_4, msg_to_check_it_7_cnu_69_in_5, msg_to_check_it_7_cnu_70_in_0, msg_to_check_it_7_cnu_70_in_1, msg_to_check_it_7_cnu_70_in_2, msg_to_check_it_7_cnu_70_in_3, msg_to_check_it_7_cnu_70_in_4, msg_to_check_it_7_cnu_70_in_5, msg_to_check_it_7_cnu_71_in_0, msg_to_check_it_7_cnu_71_in_1, msg_to_check_it_7_cnu_71_in_2, msg_to_check_it_7_cnu_71_in_3, msg_to_check_it_7_cnu_71_in_4, msg_to_check_it_7_cnu_71_in_5, msg_to_check_it_7_cnu_72_in_0, msg_to_check_it_7_cnu_72_in_1, msg_to_check_it_7_cnu_72_in_2, msg_to_check_it_7_cnu_72_in_3, msg_to_check_it_7_cnu_72_in_4, msg_to_check_it_7_cnu_72_in_5, msg_to_check_it_7_cnu_73_in_0, msg_to_check_it_7_cnu_73_in_1, msg_to_check_it_7_cnu_73_in_2, msg_to_check_it_7_cnu_73_in_3, msg_to_check_it_7_cnu_73_in_4, msg_to_check_it_7_cnu_73_in_5, msg_to_check_it_7_cnu_74_in_0, msg_to_check_it_7_cnu_74_in_1, msg_to_check_it_7_cnu_74_in_2, msg_to_check_it_7_cnu_74_in_3, msg_to_check_it_7_cnu_74_in_4, msg_to_check_it_7_cnu_74_in_5, msg_to_check_it_7_cnu_75_in_0, msg_to_check_it_7_cnu_75_in_1, msg_to_check_it_7_cnu_75_in_2, msg_to_check_it_7_cnu_75_in_3, msg_to_check_it_7_cnu_75_in_4, msg_to_check_it_7_cnu_75_in_5, msg_to_check_it_7_cnu_76_in_0, msg_to_check_it_7_cnu_76_in_1, msg_to_check_it_7_cnu_76_in_2, msg_to_check_it_7_cnu_76_in_3, msg_to_check_it_7_cnu_76_in_4, msg_to_check_it_7_cnu_76_in_5, msg_to_check_it_7_cnu_77_in_0, msg_to_check_it_7_cnu_77_in_1, msg_to_check_it_7_cnu_77_in_2, msg_to_check_it_7_cnu_77_in_3, msg_to_check_it_7_cnu_77_in_4, msg_to_check_it_7_cnu_77_in_5, msg_to_check_it_7_cnu_78_in_0, msg_to_check_it_7_cnu_78_in_1, msg_to_check_it_7_cnu_78_in_2, msg_to_check_it_7_cnu_78_in_3, msg_to_check_it_7_cnu_78_in_4, msg_to_check_it_7_cnu_78_in_5, msg_to_check_it_7_cnu_79_in_0, msg_to_check_it_7_cnu_79_in_1, msg_to_check_it_7_cnu_79_in_2, msg_to_check_it_7_cnu_79_in_3, msg_to_check_it_7_cnu_79_in_4, msg_to_check_it_7_cnu_79_in_5, msg_to_check_it_7_cnu_80_in_0, msg_to_check_it_7_cnu_80_in_1, msg_to_check_it_7_cnu_80_in_2, msg_to_check_it_7_cnu_80_in_3, msg_to_check_it_7_cnu_80_in_4, msg_to_check_it_7_cnu_80_in_5, msg_to_check_it_7_cnu_81_in_0, msg_to_check_it_7_cnu_81_in_1, msg_to_check_it_7_cnu_81_in_2, msg_to_check_it_7_cnu_81_in_3, msg_to_check_it_7_cnu_81_in_4, msg_to_check_it_7_cnu_81_in_5, msg_to_check_it_7_cnu_82_in_0, msg_to_check_it_7_cnu_82_in_1, msg_to_check_it_7_cnu_82_in_2, msg_to_check_it_7_cnu_82_in_3, msg_to_check_it_7_cnu_82_in_4, msg_to_check_it_7_cnu_82_in_5, msg_to_check_it_7_cnu_83_in_0, msg_to_check_it_7_cnu_83_in_1, msg_to_check_it_7_cnu_83_in_2, msg_to_check_it_7_cnu_83_in_3, msg_to_check_it_7_cnu_83_in_4, msg_to_check_it_7_cnu_83_in_5, msg_to_check_it_7_cnu_84_in_0, msg_to_check_it_7_cnu_84_in_1, msg_to_check_it_7_cnu_84_in_2, msg_to_check_it_7_cnu_84_in_3, msg_to_check_it_7_cnu_84_in_4, msg_to_check_it_7_cnu_84_in_5, msg_to_check_it_7_cnu_85_in_0, msg_to_check_it_7_cnu_85_in_1, msg_to_check_it_7_cnu_85_in_2, msg_to_check_it_7_cnu_85_in_3, msg_to_check_it_7_cnu_85_in_4, msg_to_check_it_7_cnu_85_in_5, msg_to_check_it_7_cnu_86_in_0, msg_to_check_it_7_cnu_86_in_1, msg_to_check_it_7_cnu_86_in_2, msg_to_check_it_7_cnu_86_in_3, msg_to_check_it_7_cnu_86_in_4, msg_to_check_it_7_cnu_86_in_5, msg_to_check_it_7_cnu_87_in_0, msg_to_check_it_7_cnu_87_in_1, msg_to_check_it_7_cnu_87_in_2, msg_to_check_it_7_cnu_87_in_3, msg_to_check_it_7_cnu_87_in_4, msg_to_check_it_7_cnu_87_in_5, msg_to_check_it_7_cnu_88_in_0, msg_to_check_it_7_cnu_88_in_1, msg_to_check_it_7_cnu_88_in_2, msg_to_check_it_7_cnu_88_in_3, msg_to_check_it_7_cnu_88_in_4, msg_to_check_it_7_cnu_88_in_5, msg_to_check_it_7_cnu_89_in_0, msg_to_check_it_7_cnu_89_in_1, msg_to_check_it_7_cnu_89_in_2, msg_to_check_it_7_cnu_89_in_3, msg_to_check_it_7_cnu_89_in_4, msg_to_check_it_7_cnu_89_in_5, msg_to_check_it_7_cnu_90_in_0, msg_to_check_it_7_cnu_90_in_1, msg_to_check_it_7_cnu_90_in_2, msg_to_check_it_7_cnu_90_in_3, msg_to_check_it_7_cnu_90_in_4, msg_to_check_it_7_cnu_90_in_5, msg_to_check_it_7_cnu_91_in_0, msg_to_check_it_7_cnu_91_in_1, msg_to_check_it_7_cnu_91_in_2, msg_to_check_it_7_cnu_91_in_3, msg_to_check_it_7_cnu_91_in_4, msg_to_check_it_7_cnu_91_in_5, msg_to_check_it_7_cnu_92_in_0, msg_to_check_it_7_cnu_92_in_1, msg_to_check_it_7_cnu_92_in_2, msg_to_check_it_7_cnu_92_in_3, msg_to_check_it_7_cnu_92_in_4, msg_to_check_it_7_cnu_92_in_5, msg_to_check_it_7_cnu_93_in_0, msg_to_check_it_7_cnu_93_in_1, msg_to_check_it_7_cnu_93_in_2, msg_to_check_it_7_cnu_93_in_3, msg_to_check_it_7_cnu_93_in_4, msg_to_check_it_7_cnu_93_in_5, msg_to_check_it_7_cnu_94_in_0, msg_to_check_it_7_cnu_94_in_1, msg_to_check_it_7_cnu_94_in_2, msg_to_check_it_7_cnu_94_in_3, msg_to_check_it_7_cnu_94_in_4, msg_to_check_it_7_cnu_94_in_5, msg_to_check_it_7_cnu_95_in_0, msg_to_check_it_7_cnu_95_in_1, msg_to_check_it_7_cnu_95_in_2, msg_to_check_it_7_cnu_95_in_3, msg_to_check_it_7_cnu_95_in_4, msg_to_check_it_7_cnu_95_in_5, msg_to_check_it_7_cnu_96_in_0, msg_to_check_it_7_cnu_96_in_1, msg_to_check_it_7_cnu_96_in_2, msg_to_check_it_7_cnu_96_in_3, msg_to_check_it_7_cnu_96_in_4, msg_to_check_it_7_cnu_96_in_5, msg_to_check_it_7_cnu_97_in_0, msg_to_check_it_7_cnu_97_in_1, msg_to_check_it_7_cnu_97_in_2, msg_to_check_it_7_cnu_97_in_3, msg_to_check_it_7_cnu_97_in_4, msg_to_check_it_7_cnu_97_in_5, msg_to_check_it_7_cnu_98_in_0, msg_to_check_it_7_cnu_98_in_1, msg_to_check_it_7_cnu_98_in_2, msg_to_check_it_7_cnu_98_in_3, msg_to_check_it_7_cnu_98_in_4, msg_to_check_it_7_cnu_98_in_5, msg_to_check_it_8_cnu_0_in_0, msg_to_check_it_8_cnu_0_in_1, msg_to_check_it_8_cnu_0_in_2, msg_to_check_it_8_cnu_0_in_3, msg_to_check_it_8_cnu_0_in_4, msg_to_check_it_8_cnu_0_in_5, msg_to_check_it_8_cnu_1_in_0, msg_to_check_it_8_cnu_1_in_1, msg_to_check_it_8_cnu_1_in_2, msg_to_check_it_8_cnu_1_in_3, msg_to_check_it_8_cnu_1_in_4, msg_to_check_it_8_cnu_1_in_5, msg_to_check_it_8_cnu_2_in_0, msg_to_check_it_8_cnu_2_in_1, msg_to_check_it_8_cnu_2_in_2, msg_to_check_it_8_cnu_2_in_3, msg_to_check_it_8_cnu_2_in_4, msg_to_check_it_8_cnu_2_in_5, msg_to_check_it_8_cnu_3_in_0, msg_to_check_it_8_cnu_3_in_1, msg_to_check_it_8_cnu_3_in_2, msg_to_check_it_8_cnu_3_in_3, msg_to_check_it_8_cnu_3_in_4, msg_to_check_it_8_cnu_3_in_5, msg_to_check_it_8_cnu_4_in_0, msg_to_check_it_8_cnu_4_in_1, msg_to_check_it_8_cnu_4_in_2, msg_to_check_it_8_cnu_4_in_3, msg_to_check_it_8_cnu_4_in_4, msg_to_check_it_8_cnu_4_in_5, msg_to_check_it_8_cnu_5_in_0, msg_to_check_it_8_cnu_5_in_1, msg_to_check_it_8_cnu_5_in_2, msg_to_check_it_8_cnu_5_in_3, msg_to_check_it_8_cnu_5_in_4, msg_to_check_it_8_cnu_5_in_5, msg_to_check_it_8_cnu_6_in_0, msg_to_check_it_8_cnu_6_in_1, msg_to_check_it_8_cnu_6_in_2, msg_to_check_it_8_cnu_6_in_3, msg_to_check_it_8_cnu_6_in_4, msg_to_check_it_8_cnu_6_in_5, msg_to_check_it_8_cnu_7_in_0, msg_to_check_it_8_cnu_7_in_1, msg_to_check_it_8_cnu_7_in_2, msg_to_check_it_8_cnu_7_in_3, msg_to_check_it_8_cnu_7_in_4, msg_to_check_it_8_cnu_7_in_5, msg_to_check_it_8_cnu_8_in_0, msg_to_check_it_8_cnu_8_in_1, msg_to_check_it_8_cnu_8_in_2, msg_to_check_it_8_cnu_8_in_3, msg_to_check_it_8_cnu_8_in_4, msg_to_check_it_8_cnu_8_in_5, msg_to_check_it_8_cnu_9_in_0, msg_to_check_it_8_cnu_9_in_1, msg_to_check_it_8_cnu_9_in_2, msg_to_check_it_8_cnu_9_in_3, msg_to_check_it_8_cnu_9_in_4, msg_to_check_it_8_cnu_9_in_5, msg_to_check_it_8_cnu_10_in_0, msg_to_check_it_8_cnu_10_in_1, msg_to_check_it_8_cnu_10_in_2, msg_to_check_it_8_cnu_10_in_3, msg_to_check_it_8_cnu_10_in_4, msg_to_check_it_8_cnu_10_in_5, msg_to_check_it_8_cnu_11_in_0, msg_to_check_it_8_cnu_11_in_1, msg_to_check_it_8_cnu_11_in_2, msg_to_check_it_8_cnu_11_in_3, msg_to_check_it_8_cnu_11_in_4, msg_to_check_it_8_cnu_11_in_5, msg_to_check_it_8_cnu_12_in_0, msg_to_check_it_8_cnu_12_in_1, msg_to_check_it_8_cnu_12_in_2, msg_to_check_it_8_cnu_12_in_3, msg_to_check_it_8_cnu_12_in_4, msg_to_check_it_8_cnu_12_in_5, msg_to_check_it_8_cnu_13_in_0, msg_to_check_it_8_cnu_13_in_1, msg_to_check_it_8_cnu_13_in_2, msg_to_check_it_8_cnu_13_in_3, msg_to_check_it_8_cnu_13_in_4, msg_to_check_it_8_cnu_13_in_5, msg_to_check_it_8_cnu_14_in_0, msg_to_check_it_8_cnu_14_in_1, msg_to_check_it_8_cnu_14_in_2, msg_to_check_it_8_cnu_14_in_3, msg_to_check_it_8_cnu_14_in_4, msg_to_check_it_8_cnu_14_in_5, msg_to_check_it_8_cnu_15_in_0, msg_to_check_it_8_cnu_15_in_1, msg_to_check_it_8_cnu_15_in_2, msg_to_check_it_8_cnu_15_in_3, msg_to_check_it_8_cnu_15_in_4, msg_to_check_it_8_cnu_15_in_5, msg_to_check_it_8_cnu_16_in_0, msg_to_check_it_8_cnu_16_in_1, msg_to_check_it_8_cnu_16_in_2, msg_to_check_it_8_cnu_16_in_3, msg_to_check_it_8_cnu_16_in_4, msg_to_check_it_8_cnu_16_in_5, msg_to_check_it_8_cnu_17_in_0, msg_to_check_it_8_cnu_17_in_1, msg_to_check_it_8_cnu_17_in_2, msg_to_check_it_8_cnu_17_in_3, msg_to_check_it_8_cnu_17_in_4, msg_to_check_it_8_cnu_17_in_5, msg_to_check_it_8_cnu_18_in_0, msg_to_check_it_8_cnu_18_in_1, msg_to_check_it_8_cnu_18_in_2, msg_to_check_it_8_cnu_18_in_3, msg_to_check_it_8_cnu_18_in_4, msg_to_check_it_8_cnu_18_in_5, msg_to_check_it_8_cnu_19_in_0, msg_to_check_it_8_cnu_19_in_1, msg_to_check_it_8_cnu_19_in_2, msg_to_check_it_8_cnu_19_in_3, msg_to_check_it_8_cnu_19_in_4, msg_to_check_it_8_cnu_19_in_5, msg_to_check_it_8_cnu_20_in_0, msg_to_check_it_8_cnu_20_in_1, msg_to_check_it_8_cnu_20_in_2, msg_to_check_it_8_cnu_20_in_3, msg_to_check_it_8_cnu_20_in_4, msg_to_check_it_8_cnu_20_in_5, msg_to_check_it_8_cnu_21_in_0, msg_to_check_it_8_cnu_21_in_1, msg_to_check_it_8_cnu_21_in_2, msg_to_check_it_8_cnu_21_in_3, msg_to_check_it_8_cnu_21_in_4, msg_to_check_it_8_cnu_21_in_5, msg_to_check_it_8_cnu_22_in_0, msg_to_check_it_8_cnu_22_in_1, msg_to_check_it_8_cnu_22_in_2, msg_to_check_it_8_cnu_22_in_3, msg_to_check_it_8_cnu_22_in_4, msg_to_check_it_8_cnu_22_in_5, msg_to_check_it_8_cnu_23_in_0, msg_to_check_it_8_cnu_23_in_1, msg_to_check_it_8_cnu_23_in_2, msg_to_check_it_8_cnu_23_in_3, msg_to_check_it_8_cnu_23_in_4, msg_to_check_it_8_cnu_23_in_5, msg_to_check_it_8_cnu_24_in_0, msg_to_check_it_8_cnu_24_in_1, msg_to_check_it_8_cnu_24_in_2, msg_to_check_it_8_cnu_24_in_3, msg_to_check_it_8_cnu_24_in_4, msg_to_check_it_8_cnu_24_in_5, msg_to_check_it_8_cnu_25_in_0, msg_to_check_it_8_cnu_25_in_1, msg_to_check_it_8_cnu_25_in_2, msg_to_check_it_8_cnu_25_in_3, msg_to_check_it_8_cnu_25_in_4, msg_to_check_it_8_cnu_25_in_5, msg_to_check_it_8_cnu_26_in_0, msg_to_check_it_8_cnu_26_in_1, msg_to_check_it_8_cnu_26_in_2, msg_to_check_it_8_cnu_26_in_3, msg_to_check_it_8_cnu_26_in_4, msg_to_check_it_8_cnu_26_in_5, msg_to_check_it_8_cnu_27_in_0, msg_to_check_it_8_cnu_27_in_1, msg_to_check_it_8_cnu_27_in_2, msg_to_check_it_8_cnu_27_in_3, msg_to_check_it_8_cnu_27_in_4, msg_to_check_it_8_cnu_27_in_5, msg_to_check_it_8_cnu_28_in_0, msg_to_check_it_8_cnu_28_in_1, msg_to_check_it_8_cnu_28_in_2, msg_to_check_it_8_cnu_28_in_3, msg_to_check_it_8_cnu_28_in_4, msg_to_check_it_8_cnu_28_in_5, msg_to_check_it_8_cnu_29_in_0, msg_to_check_it_8_cnu_29_in_1, msg_to_check_it_8_cnu_29_in_2, msg_to_check_it_8_cnu_29_in_3, msg_to_check_it_8_cnu_29_in_4, msg_to_check_it_8_cnu_29_in_5, msg_to_check_it_8_cnu_30_in_0, msg_to_check_it_8_cnu_30_in_1, msg_to_check_it_8_cnu_30_in_2, msg_to_check_it_8_cnu_30_in_3, msg_to_check_it_8_cnu_30_in_4, msg_to_check_it_8_cnu_30_in_5, msg_to_check_it_8_cnu_31_in_0, msg_to_check_it_8_cnu_31_in_1, msg_to_check_it_8_cnu_31_in_2, msg_to_check_it_8_cnu_31_in_3, msg_to_check_it_8_cnu_31_in_4, msg_to_check_it_8_cnu_31_in_5, msg_to_check_it_8_cnu_32_in_0, msg_to_check_it_8_cnu_32_in_1, msg_to_check_it_8_cnu_32_in_2, msg_to_check_it_8_cnu_32_in_3, msg_to_check_it_8_cnu_32_in_4, msg_to_check_it_8_cnu_32_in_5, msg_to_check_it_8_cnu_33_in_0, msg_to_check_it_8_cnu_33_in_1, msg_to_check_it_8_cnu_33_in_2, msg_to_check_it_8_cnu_33_in_3, msg_to_check_it_8_cnu_33_in_4, msg_to_check_it_8_cnu_33_in_5, msg_to_check_it_8_cnu_34_in_0, msg_to_check_it_8_cnu_34_in_1, msg_to_check_it_8_cnu_34_in_2, msg_to_check_it_8_cnu_34_in_3, msg_to_check_it_8_cnu_34_in_4, msg_to_check_it_8_cnu_34_in_5, msg_to_check_it_8_cnu_35_in_0, msg_to_check_it_8_cnu_35_in_1, msg_to_check_it_8_cnu_35_in_2, msg_to_check_it_8_cnu_35_in_3, msg_to_check_it_8_cnu_35_in_4, msg_to_check_it_8_cnu_35_in_5, msg_to_check_it_8_cnu_36_in_0, msg_to_check_it_8_cnu_36_in_1, msg_to_check_it_8_cnu_36_in_2, msg_to_check_it_8_cnu_36_in_3, msg_to_check_it_8_cnu_36_in_4, msg_to_check_it_8_cnu_36_in_5, msg_to_check_it_8_cnu_37_in_0, msg_to_check_it_8_cnu_37_in_1, msg_to_check_it_8_cnu_37_in_2, msg_to_check_it_8_cnu_37_in_3, msg_to_check_it_8_cnu_37_in_4, msg_to_check_it_8_cnu_37_in_5, msg_to_check_it_8_cnu_38_in_0, msg_to_check_it_8_cnu_38_in_1, msg_to_check_it_8_cnu_38_in_2, msg_to_check_it_8_cnu_38_in_3, msg_to_check_it_8_cnu_38_in_4, msg_to_check_it_8_cnu_38_in_5, msg_to_check_it_8_cnu_39_in_0, msg_to_check_it_8_cnu_39_in_1, msg_to_check_it_8_cnu_39_in_2, msg_to_check_it_8_cnu_39_in_3, msg_to_check_it_8_cnu_39_in_4, msg_to_check_it_8_cnu_39_in_5, msg_to_check_it_8_cnu_40_in_0, msg_to_check_it_8_cnu_40_in_1, msg_to_check_it_8_cnu_40_in_2, msg_to_check_it_8_cnu_40_in_3, msg_to_check_it_8_cnu_40_in_4, msg_to_check_it_8_cnu_40_in_5, msg_to_check_it_8_cnu_41_in_0, msg_to_check_it_8_cnu_41_in_1, msg_to_check_it_8_cnu_41_in_2, msg_to_check_it_8_cnu_41_in_3, msg_to_check_it_8_cnu_41_in_4, msg_to_check_it_8_cnu_41_in_5, msg_to_check_it_8_cnu_42_in_0, msg_to_check_it_8_cnu_42_in_1, msg_to_check_it_8_cnu_42_in_2, msg_to_check_it_8_cnu_42_in_3, msg_to_check_it_8_cnu_42_in_4, msg_to_check_it_8_cnu_42_in_5, msg_to_check_it_8_cnu_43_in_0, msg_to_check_it_8_cnu_43_in_1, msg_to_check_it_8_cnu_43_in_2, msg_to_check_it_8_cnu_43_in_3, msg_to_check_it_8_cnu_43_in_4, msg_to_check_it_8_cnu_43_in_5, msg_to_check_it_8_cnu_44_in_0, msg_to_check_it_8_cnu_44_in_1, msg_to_check_it_8_cnu_44_in_2, msg_to_check_it_8_cnu_44_in_3, msg_to_check_it_8_cnu_44_in_4, msg_to_check_it_8_cnu_44_in_5, msg_to_check_it_8_cnu_45_in_0, msg_to_check_it_8_cnu_45_in_1, msg_to_check_it_8_cnu_45_in_2, msg_to_check_it_8_cnu_45_in_3, msg_to_check_it_8_cnu_45_in_4, msg_to_check_it_8_cnu_45_in_5, msg_to_check_it_8_cnu_46_in_0, msg_to_check_it_8_cnu_46_in_1, msg_to_check_it_8_cnu_46_in_2, msg_to_check_it_8_cnu_46_in_3, msg_to_check_it_8_cnu_46_in_4, msg_to_check_it_8_cnu_46_in_5, msg_to_check_it_8_cnu_47_in_0, msg_to_check_it_8_cnu_47_in_1, msg_to_check_it_8_cnu_47_in_2, msg_to_check_it_8_cnu_47_in_3, msg_to_check_it_8_cnu_47_in_4, msg_to_check_it_8_cnu_47_in_5, msg_to_check_it_8_cnu_48_in_0, msg_to_check_it_8_cnu_48_in_1, msg_to_check_it_8_cnu_48_in_2, msg_to_check_it_8_cnu_48_in_3, msg_to_check_it_8_cnu_48_in_4, msg_to_check_it_8_cnu_48_in_5, msg_to_check_it_8_cnu_49_in_0, msg_to_check_it_8_cnu_49_in_1, msg_to_check_it_8_cnu_49_in_2, msg_to_check_it_8_cnu_49_in_3, msg_to_check_it_8_cnu_49_in_4, msg_to_check_it_8_cnu_49_in_5, msg_to_check_it_8_cnu_50_in_0, msg_to_check_it_8_cnu_50_in_1, msg_to_check_it_8_cnu_50_in_2, msg_to_check_it_8_cnu_50_in_3, msg_to_check_it_8_cnu_50_in_4, msg_to_check_it_8_cnu_50_in_5, msg_to_check_it_8_cnu_51_in_0, msg_to_check_it_8_cnu_51_in_1, msg_to_check_it_8_cnu_51_in_2, msg_to_check_it_8_cnu_51_in_3, msg_to_check_it_8_cnu_51_in_4, msg_to_check_it_8_cnu_51_in_5, msg_to_check_it_8_cnu_52_in_0, msg_to_check_it_8_cnu_52_in_1, msg_to_check_it_8_cnu_52_in_2, msg_to_check_it_8_cnu_52_in_3, msg_to_check_it_8_cnu_52_in_4, msg_to_check_it_8_cnu_52_in_5, msg_to_check_it_8_cnu_53_in_0, msg_to_check_it_8_cnu_53_in_1, msg_to_check_it_8_cnu_53_in_2, msg_to_check_it_8_cnu_53_in_3, msg_to_check_it_8_cnu_53_in_4, msg_to_check_it_8_cnu_53_in_5, msg_to_check_it_8_cnu_54_in_0, msg_to_check_it_8_cnu_54_in_1, msg_to_check_it_8_cnu_54_in_2, msg_to_check_it_8_cnu_54_in_3, msg_to_check_it_8_cnu_54_in_4, msg_to_check_it_8_cnu_54_in_5, msg_to_check_it_8_cnu_55_in_0, msg_to_check_it_8_cnu_55_in_1, msg_to_check_it_8_cnu_55_in_2, msg_to_check_it_8_cnu_55_in_3, msg_to_check_it_8_cnu_55_in_4, msg_to_check_it_8_cnu_55_in_5, msg_to_check_it_8_cnu_56_in_0, msg_to_check_it_8_cnu_56_in_1, msg_to_check_it_8_cnu_56_in_2, msg_to_check_it_8_cnu_56_in_3, msg_to_check_it_8_cnu_56_in_4, msg_to_check_it_8_cnu_56_in_5, msg_to_check_it_8_cnu_57_in_0, msg_to_check_it_8_cnu_57_in_1, msg_to_check_it_8_cnu_57_in_2, msg_to_check_it_8_cnu_57_in_3, msg_to_check_it_8_cnu_57_in_4, msg_to_check_it_8_cnu_57_in_5, msg_to_check_it_8_cnu_58_in_0, msg_to_check_it_8_cnu_58_in_1, msg_to_check_it_8_cnu_58_in_2, msg_to_check_it_8_cnu_58_in_3, msg_to_check_it_8_cnu_58_in_4, msg_to_check_it_8_cnu_58_in_5, msg_to_check_it_8_cnu_59_in_0, msg_to_check_it_8_cnu_59_in_1, msg_to_check_it_8_cnu_59_in_2, msg_to_check_it_8_cnu_59_in_3, msg_to_check_it_8_cnu_59_in_4, msg_to_check_it_8_cnu_59_in_5, msg_to_check_it_8_cnu_60_in_0, msg_to_check_it_8_cnu_60_in_1, msg_to_check_it_8_cnu_60_in_2, msg_to_check_it_8_cnu_60_in_3, msg_to_check_it_8_cnu_60_in_4, msg_to_check_it_8_cnu_60_in_5, msg_to_check_it_8_cnu_61_in_0, msg_to_check_it_8_cnu_61_in_1, msg_to_check_it_8_cnu_61_in_2, msg_to_check_it_8_cnu_61_in_3, msg_to_check_it_8_cnu_61_in_4, msg_to_check_it_8_cnu_61_in_5, msg_to_check_it_8_cnu_62_in_0, msg_to_check_it_8_cnu_62_in_1, msg_to_check_it_8_cnu_62_in_2, msg_to_check_it_8_cnu_62_in_3, msg_to_check_it_8_cnu_62_in_4, msg_to_check_it_8_cnu_62_in_5, msg_to_check_it_8_cnu_63_in_0, msg_to_check_it_8_cnu_63_in_1, msg_to_check_it_8_cnu_63_in_2, msg_to_check_it_8_cnu_63_in_3, msg_to_check_it_8_cnu_63_in_4, msg_to_check_it_8_cnu_63_in_5, msg_to_check_it_8_cnu_64_in_0, msg_to_check_it_8_cnu_64_in_1, msg_to_check_it_8_cnu_64_in_2, msg_to_check_it_8_cnu_64_in_3, msg_to_check_it_8_cnu_64_in_4, msg_to_check_it_8_cnu_64_in_5, msg_to_check_it_8_cnu_65_in_0, msg_to_check_it_8_cnu_65_in_1, msg_to_check_it_8_cnu_65_in_2, msg_to_check_it_8_cnu_65_in_3, msg_to_check_it_8_cnu_65_in_4, msg_to_check_it_8_cnu_65_in_5, msg_to_check_it_8_cnu_66_in_0, msg_to_check_it_8_cnu_66_in_1, msg_to_check_it_8_cnu_66_in_2, msg_to_check_it_8_cnu_66_in_3, msg_to_check_it_8_cnu_66_in_4, msg_to_check_it_8_cnu_66_in_5, msg_to_check_it_8_cnu_67_in_0, msg_to_check_it_8_cnu_67_in_1, msg_to_check_it_8_cnu_67_in_2, msg_to_check_it_8_cnu_67_in_3, msg_to_check_it_8_cnu_67_in_4, msg_to_check_it_8_cnu_67_in_5, msg_to_check_it_8_cnu_68_in_0, msg_to_check_it_8_cnu_68_in_1, msg_to_check_it_8_cnu_68_in_2, msg_to_check_it_8_cnu_68_in_3, msg_to_check_it_8_cnu_68_in_4, msg_to_check_it_8_cnu_68_in_5, msg_to_check_it_8_cnu_69_in_0, msg_to_check_it_8_cnu_69_in_1, msg_to_check_it_8_cnu_69_in_2, msg_to_check_it_8_cnu_69_in_3, msg_to_check_it_8_cnu_69_in_4, msg_to_check_it_8_cnu_69_in_5, msg_to_check_it_8_cnu_70_in_0, msg_to_check_it_8_cnu_70_in_1, msg_to_check_it_8_cnu_70_in_2, msg_to_check_it_8_cnu_70_in_3, msg_to_check_it_8_cnu_70_in_4, msg_to_check_it_8_cnu_70_in_5, msg_to_check_it_8_cnu_71_in_0, msg_to_check_it_8_cnu_71_in_1, msg_to_check_it_8_cnu_71_in_2, msg_to_check_it_8_cnu_71_in_3, msg_to_check_it_8_cnu_71_in_4, msg_to_check_it_8_cnu_71_in_5, msg_to_check_it_8_cnu_72_in_0, msg_to_check_it_8_cnu_72_in_1, msg_to_check_it_8_cnu_72_in_2, msg_to_check_it_8_cnu_72_in_3, msg_to_check_it_8_cnu_72_in_4, msg_to_check_it_8_cnu_72_in_5, msg_to_check_it_8_cnu_73_in_0, msg_to_check_it_8_cnu_73_in_1, msg_to_check_it_8_cnu_73_in_2, msg_to_check_it_8_cnu_73_in_3, msg_to_check_it_8_cnu_73_in_4, msg_to_check_it_8_cnu_73_in_5, msg_to_check_it_8_cnu_74_in_0, msg_to_check_it_8_cnu_74_in_1, msg_to_check_it_8_cnu_74_in_2, msg_to_check_it_8_cnu_74_in_3, msg_to_check_it_8_cnu_74_in_4, msg_to_check_it_8_cnu_74_in_5, msg_to_check_it_8_cnu_75_in_0, msg_to_check_it_8_cnu_75_in_1, msg_to_check_it_8_cnu_75_in_2, msg_to_check_it_8_cnu_75_in_3, msg_to_check_it_8_cnu_75_in_4, msg_to_check_it_8_cnu_75_in_5, msg_to_check_it_8_cnu_76_in_0, msg_to_check_it_8_cnu_76_in_1, msg_to_check_it_8_cnu_76_in_2, msg_to_check_it_8_cnu_76_in_3, msg_to_check_it_8_cnu_76_in_4, msg_to_check_it_8_cnu_76_in_5, msg_to_check_it_8_cnu_77_in_0, msg_to_check_it_8_cnu_77_in_1, msg_to_check_it_8_cnu_77_in_2, msg_to_check_it_8_cnu_77_in_3, msg_to_check_it_8_cnu_77_in_4, msg_to_check_it_8_cnu_77_in_5, msg_to_check_it_8_cnu_78_in_0, msg_to_check_it_8_cnu_78_in_1, msg_to_check_it_8_cnu_78_in_2, msg_to_check_it_8_cnu_78_in_3, msg_to_check_it_8_cnu_78_in_4, msg_to_check_it_8_cnu_78_in_5, msg_to_check_it_8_cnu_79_in_0, msg_to_check_it_8_cnu_79_in_1, msg_to_check_it_8_cnu_79_in_2, msg_to_check_it_8_cnu_79_in_3, msg_to_check_it_8_cnu_79_in_4, msg_to_check_it_8_cnu_79_in_5, msg_to_check_it_8_cnu_80_in_0, msg_to_check_it_8_cnu_80_in_1, msg_to_check_it_8_cnu_80_in_2, msg_to_check_it_8_cnu_80_in_3, msg_to_check_it_8_cnu_80_in_4, msg_to_check_it_8_cnu_80_in_5, msg_to_check_it_8_cnu_81_in_0, msg_to_check_it_8_cnu_81_in_1, msg_to_check_it_8_cnu_81_in_2, msg_to_check_it_8_cnu_81_in_3, msg_to_check_it_8_cnu_81_in_4, msg_to_check_it_8_cnu_81_in_5, msg_to_check_it_8_cnu_82_in_0, msg_to_check_it_8_cnu_82_in_1, msg_to_check_it_8_cnu_82_in_2, msg_to_check_it_8_cnu_82_in_3, msg_to_check_it_8_cnu_82_in_4, msg_to_check_it_8_cnu_82_in_5, msg_to_check_it_8_cnu_83_in_0, msg_to_check_it_8_cnu_83_in_1, msg_to_check_it_8_cnu_83_in_2, msg_to_check_it_8_cnu_83_in_3, msg_to_check_it_8_cnu_83_in_4, msg_to_check_it_8_cnu_83_in_5, msg_to_check_it_8_cnu_84_in_0, msg_to_check_it_8_cnu_84_in_1, msg_to_check_it_8_cnu_84_in_2, msg_to_check_it_8_cnu_84_in_3, msg_to_check_it_8_cnu_84_in_4, msg_to_check_it_8_cnu_84_in_5, msg_to_check_it_8_cnu_85_in_0, msg_to_check_it_8_cnu_85_in_1, msg_to_check_it_8_cnu_85_in_2, msg_to_check_it_8_cnu_85_in_3, msg_to_check_it_8_cnu_85_in_4, msg_to_check_it_8_cnu_85_in_5, msg_to_check_it_8_cnu_86_in_0, msg_to_check_it_8_cnu_86_in_1, msg_to_check_it_8_cnu_86_in_2, msg_to_check_it_8_cnu_86_in_3, msg_to_check_it_8_cnu_86_in_4, msg_to_check_it_8_cnu_86_in_5, msg_to_check_it_8_cnu_87_in_0, msg_to_check_it_8_cnu_87_in_1, msg_to_check_it_8_cnu_87_in_2, msg_to_check_it_8_cnu_87_in_3, msg_to_check_it_8_cnu_87_in_4, msg_to_check_it_8_cnu_87_in_5, msg_to_check_it_8_cnu_88_in_0, msg_to_check_it_8_cnu_88_in_1, msg_to_check_it_8_cnu_88_in_2, msg_to_check_it_8_cnu_88_in_3, msg_to_check_it_8_cnu_88_in_4, msg_to_check_it_8_cnu_88_in_5, msg_to_check_it_8_cnu_89_in_0, msg_to_check_it_8_cnu_89_in_1, msg_to_check_it_8_cnu_89_in_2, msg_to_check_it_8_cnu_89_in_3, msg_to_check_it_8_cnu_89_in_4, msg_to_check_it_8_cnu_89_in_5, msg_to_check_it_8_cnu_90_in_0, msg_to_check_it_8_cnu_90_in_1, msg_to_check_it_8_cnu_90_in_2, msg_to_check_it_8_cnu_90_in_3, msg_to_check_it_8_cnu_90_in_4, msg_to_check_it_8_cnu_90_in_5, msg_to_check_it_8_cnu_91_in_0, msg_to_check_it_8_cnu_91_in_1, msg_to_check_it_8_cnu_91_in_2, msg_to_check_it_8_cnu_91_in_3, msg_to_check_it_8_cnu_91_in_4, msg_to_check_it_8_cnu_91_in_5, msg_to_check_it_8_cnu_92_in_0, msg_to_check_it_8_cnu_92_in_1, msg_to_check_it_8_cnu_92_in_2, msg_to_check_it_8_cnu_92_in_3, msg_to_check_it_8_cnu_92_in_4, msg_to_check_it_8_cnu_92_in_5, msg_to_check_it_8_cnu_93_in_0, msg_to_check_it_8_cnu_93_in_1, msg_to_check_it_8_cnu_93_in_2, msg_to_check_it_8_cnu_93_in_3, msg_to_check_it_8_cnu_93_in_4, msg_to_check_it_8_cnu_93_in_5, msg_to_check_it_8_cnu_94_in_0, msg_to_check_it_8_cnu_94_in_1, msg_to_check_it_8_cnu_94_in_2, msg_to_check_it_8_cnu_94_in_3, msg_to_check_it_8_cnu_94_in_4, msg_to_check_it_8_cnu_94_in_5, msg_to_check_it_8_cnu_95_in_0, msg_to_check_it_8_cnu_95_in_1, msg_to_check_it_8_cnu_95_in_2, msg_to_check_it_8_cnu_95_in_3, msg_to_check_it_8_cnu_95_in_4, msg_to_check_it_8_cnu_95_in_5, msg_to_check_it_8_cnu_96_in_0, msg_to_check_it_8_cnu_96_in_1, msg_to_check_it_8_cnu_96_in_2, msg_to_check_it_8_cnu_96_in_3, msg_to_check_it_8_cnu_96_in_4, msg_to_check_it_8_cnu_96_in_5, msg_to_check_it_8_cnu_97_in_0, msg_to_check_it_8_cnu_97_in_1, msg_to_check_it_8_cnu_97_in_2, msg_to_check_it_8_cnu_97_in_3, msg_to_check_it_8_cnu_97_in_4, msg_to_check_it_8_cnu_97_in_5, msg_to_check_it_8_cnu_98_in_0, msg_to_check_it_8_cnu_98_in_1, msg_to_check_it_8_cnu_98_in_2, msg_to_check_it_8_cnu_98_in_3, msg_to_check_it_8_cnu_98_in_4, msg_to_check_it_8_cnu_98_in_5, msg_to_check_it_9_cnu_0_in_0, msg_to_check_it_9_cnu_0_in_1, msg_to_check_it_9_cnu_0_in_2, msg_to_check_it_9_cnu_0_in_3, msg_to_check_it_9_cnu_0_in_4, msg_to_check_it_9_cnu_0_in_5, msg_to_check_it_9_cnu_1_in_0, msg_to_check_it_9_cnu_1_in_1, msg_to_check_it_9_cnu_1_in_2, msg_to_check_it_9_cnu_1_in_3, msg_to_check_it_9_cnu_1_in_4, msg_to_check_it_9_cnu_1_in_5, msg_to_check_it_9_cnu_2_in_0, msg_to_check_it_9_cnu_2_in_1, msg_to_check_it_9_cnu_2_in_2, msg_to_check_it_9_cnu_2_in_3, msg_to_check_it_9_cnu_2_in_4, msg_to_check_it_9_cnu_2_in_5, msg_to_check_it_9_cnu_3_in_0, msg_to_check_it_9_cnu_3_in_1, msg_to_check_it_9_cnu_3_in_2, msg_to_check_it_9_cnu_3_in_3, msg_to_check_it_9_cnu_3_in_4, msg_to_check_it_9_cnu_3_in_5, msg_to_check_it_9_cnu_4_in_0, msg_to_check_it_9_cnu_4_in_1, msg_to_check_it_9_cnu_4_in_2, msg_to_check_it_9_cnu_4_in_3, msg_to_check_it_9_cnu_4_in_4, msg_to_check_it_9_cnu_4_in_5, msg_to_check_it_9_cnu_5_in_0, msg_to_check_it_9_cnu_5_in_1, msg_to_check_it_9_cnu_5_in_2, msg_to_check_it_9_cnu_5_in_3, msg_to_check_it_9_cnu_5_in_4, msg_to_check_it_9_cnu_5_in_5, msg_to_check_it_9_cnu_6_in_0, msg_to_check_it_9_cnu_6_in_1, msg_to_check_it_9_cnu_6_in_2, msg_to_check_it_9_cnu_6_in_3, msg_to_check_it_9_cnu_6_in_4, msg_to_check_it_9_cnu_6_in_5, msg_to_check_it_9_cnu_7_in_0, msg_to_check_it_9_cnu_7_in_1, msg_to_check_it_9_cnu_7_in_2, msg_to_check_it_9_cnu_7_in_3, msg_to_check_it_9_cnu_7_in_4, msg_to_check_it_9_cnu_7_in_5, msg_to_check_it_9_cnu_8_in_0, msg_to_check_it_9_cnu_8_in_1, msg_to_check_it_9_cnu_8_in_2, msg_to_check_it_9_cnu_8_in_3, msg_to_check_it_9_cnu_8_in_4, msg_to_check_it_9_cnu_8_in_5, msg_to_check_it_9_cnu_9_in_0, msg_to_check_it_9_cnu_9_in_1, msg_to_check_it_9_cnu_9_in_2, msg_to_check_it_9_cnu_9_in_3, msg_to_check_it_9_cnu_9_in_4, msg_to_check_it_9_cnu_9_in_5, msg_to_check_it_9_cnu_10_in_0, msg_to_check_it_9_cnu_10_in_1, msg_to_check_it_9_cnu_10_in_2, msg_to_check_it_9_cnu_10_in_3, msg_to_check_it_9_cnu_10_in_4, msg_to_check_it_9_cnu_10_in_5, msg_to_check_it_9_cnu_11_in_0, msg_to_check_it_9_cnu_11_in_1, msg_to_check_it_9_cnu_11_in_2, msg_to_check_it_9_cnu_11_in_3, msg_to_check_it_9_cnu_11_in_4, msg_to_check_it_9_cnu_11_in_5, msg_to_check_it_9_cnu_12_in_0, msg_to_check_it_9_cnu_12_in_1, msg_to_check_it_9_cnu_12_in_2, msg_to_check_it_9_cnu_12_in_3, msg_to_check_it_9_cnu_12_in_4, msg_to_check_it_9_cnu_12_in_5, msg_to_check_it_9_cnu_13_in_0, msg_to_check_it_9_cnu_13_in_1, msg_to_check_it_9_cnu_13_in_2, msg_to_check_it_9_cnu_13_in_3, msg_to_check_it_9_cnu_13_in_4, msg_to_check_it_9_cnu_13_in_5, msg_to_check_it_9_cnu_14_in_0, msg_to_check_it_9_cnu_14_in_1, msg_to_check_it_9_cnu_14_in_2, msg_to_check_it_9_cnu_14_in_3, msg_to_check_it_9_cnu_14_in_4, msg_to_check_it_9_cnu_14_in_5, msg_to_check_it_9_cnu_15_in_0, msg_to_check_it_9_cnu_15_in_1, msg_to_check_it_9_cnu_15_in_2, msg_to_check_it_9_cnu_15_in_3, msg_to_check_it_9_cnu_15_in_4, msg_to_check_it_9_cnu_15_in_5, msg_to_check_it_9_cnu_16_in_0, msg_to_check_it_9_cnu_16_in_1, msg_to_check_it_9_cnu_16_in_2, msg_to_check_it_9_cnu_16_in_3, msg_to_check_it_9_cnu_16_in_4, msg_to_check_it_9_cnu_16_in_5, msg_to_check_it_9_cnu_17_in_0, msg_to_check_it_9_cnu_17_in_1, msg_to_check_it_9_cnu_17_in_2, msg_to_check_it_9_cnu_17_in_3, msg_to_check_it_9_cnu_17_in_4, msg_to_check_it_9_cnu_17_in_5, msg_to_check_it_9_cnu_18_in_0, msg_to_check_it_9_cnu_18_in_1, msg_to_check_it_9_cnu_18_in_2, msg_to_check_it_9_cnu_18_in_3, msg_to_check_it_9_cnu_18_in_4, msg_to_check_it_9_cnu_18_in_5, msg_to_check_it_9_cnu_19_in_0, msg_to_check_it_9_cnu_19_in_1, msg_to_check_it_9_cnu_19_in_2, msg_to_check_it_9_cnu_19_in_3, msg_to_check_it_9_cnu_19_in_4, msg_to_check_it_9_cnu_19_in_5, msg_to_check_it_9_cnu_20_in_0, msg_to_check_it_9_cnu_20_in_1, msg_to_check_it_9_cnu_20_in_2, msg_to_check_it_9_cnu_20_in_3, msg_to_check_it_9_cnu_20_in_4, msg_to_check_it_9_cnu_20_in_5, msg_to_check_it_9_cnu_21_in_0, msg_to_check_it_9_cnu_21_in_1, msg_to_check_it_9_cnu_21_in_2, msg_to_check_it_9_cnu_21_in_3, msg_to_check_it_9_cnu_21_in_4, msg_to_check_it_9_cnu_21_in_5, msg_to_check_it_9_cnu_22_in_0, msg_to_check_it_9_cnu_22_in_1, msg_to_check_it_9_cnu_22_in_2, msg_to_check_it_9_cnu_22_in_3, msg_to_check_it_9_cnu_22_in_4, msg_to_check_it_9_cnu_22_in_5, msg_to_check_it_9_cnu_23_in_0, msg_to_check_it_9_cnu_23_in_1, msg_to_check_it_9_cnu_23_in_2, msg_to_check_it_9_cnu_23_in_3, msg_to_check_it_9_cnu_23_in_4, msg_to_check_it_9_cnu_23_in_5, msg_to_check_it_9_cnu_24_in_0, msg_to_check_it_9_cnu_24_in_1, msg_to_check_it_9_cnu_24_in_2, msg_to_check_it_9_cnu_24_in_3, msg_to_check_it_9_cnu_24_in_4, msg_to_check_it_9_cnu_24_in_5, msg_to_check_it_9_cnu_25_in_0, msg_to_check_it_9_cnu_25_in_1, msg_to_check_it_9_cnu_25_in_2, msg_to_check_it_9_cnu_25_in_3, msg_to_check_it_9_cnu_25_in_4, msg_to_check_it_9_cnu_25_in_5, msg_to_check_it_9_cnu_26_in_0, msg_to_check_it_9_cnu_26_in_1, msg_to_check_it_9_cnu_26_in_2, msg_to_check_it_9_cnu_26_in_3, msg_to_check_it_9_cnu_26_in_4, msg_to_check_it_9_cnu_26_in_5, msg_to_check_it_9_cnu_27_in_0, msg_to_check_it_9_cnu_27_in_1, msg_to_check_it_9_cnu_27_in_2, msg_to_check_it_9_cnu_27_in_3, msg_to_check_it_9_cnu_27_in_4, msg_to_check_it_9_cnu_27_in_5, msg_to_check_it_9_cnu_28_in_0, msg_to_check_it_9_cnu_28_in_1, msg_to_check_it_9_cnu_28_in_2, msg_to_check_it_9_cnu_28_in_3, msg_to_check_it_9_cnu_28_in_4, msg_to_check_it_9_cnu_28_in_5, msg_to_check_it_9_cnu_29_in_0, msg_to_check_it_9_cnu_29_in_1, msg_to_check_it_9_cnu_29_in_2, msg_to_check_it_9_cnu_29_in_3, msg_to_check_it_9_cnu_29_in_4, msg_to_check_it_9_cnu_29_in_5, msg_to_check_it_9_cnu_30_in_0, msg_to_check_it_9_cnu_30_in_1, msg_to_check_it_9_cnu_30_in_2, msg_to_check_it_9_cnu_30_in_3, msg_to_check_it_9_cnu_30_in_4, msg_to_check_it_9_cnu_30_in_5, msg_to_check_it_9_cnu_31_in_0, msg_to_check_it_9_cnu_31_in_1, msg_to_check_it_9_cnu_31_in_2, msg_to_check_it_9_cnu_31_in_3, msg_to_check_it_9_cnu_31_in_4, msg_to_check_it_9_cnu_31_in_5, msg_to_check_it_9_cnu_32_in_0, msg_to_check_it_9_cnu_32_in_1, msg_to_check_it_9_cnu_32_in_2, msg_to_check_it_9_cnu_32_in_3, msg_to_check_it_9_cnu_32_in_4, msg_to_check_it_9_cnu_32_in_5, msg_to_check_it_9_cnu_33_in_0, msg_to_check_it_9_cnu_33_in_1, msg_to_check_it_9_cnu_33_in_2, msg_to_check_it_9_cnu_33_in_3, msg_to_check_it_9_cnu_33_in_4, msg_to_check_it_9_cnu_33_in_5, msg_to_check_it_9_cnu_34_in_0, msg_to_check_it_9_cnu_34_in_1, msg_to_check_it_9_cnu_34_in_2, msg_to_check_it_9_cnu_34_in_3, msg_to_check_it_9_cnu_34_in_4, msg_to_check_it_9_cnu_34_in_5, msg_to_check_it_9_cnu_35_in_0, msg_to_check_it_9_cnu_35_in_1, msg_to_check_it_9_cnu_35_in_2, msg_to_check_it_9_cnu_35_in_3, msg_to_check_it_9_cnu_35_in_4, msg_to_check_it_9_cnu_35_in_5, msg_to_check_it_9_cnu_36_in_0, msg_to_check_it_9_cnu_36_in_1, msg_to_check_it_9_cnu_36_in_2, msg_to_check_it_9_cnu_36_in_3, msg_to_check_it_9_cnu_36_in_4, msg_to_check_it_9_cnu_36_in_5, msg_to_check_it_9_cnu_37_in_0, msg_to_check_it_9_cnu_37_in_1, msg_to_check_it_9_cnu_37_in_2, msg_to_check_it_9_cnu_37_in_3, msg_to_check_it_9_cnu_37_in_4, msg_to_check_it_9_cnu_37_in_5, msg_to_check_it_9_cnu_38_in_0, msg_to_check_it_9_cnu_38_in_1, msg_to_check_it_9_cnu_38_in_2, msg_to_check_it_9_cnu_38_in_3, msg_to_check_it_9_cnu_38_in_4, msg_to_check_it_9_cnu_38_in_5, msg_to_check_it_9_cnu_39_in_0, msg_to_check_it_9_cnu_39_in_1, msg_to_check_it_9_cnu_39_in_2, msg_to_check_it_9_cnu_39_in_3, msg_to_check_it_9_cnu_39_in_4, msg_to_check_it_9_cnu_39_in_5, msg_to_check_it_9_cnu_40_in_0, msg_to_check_it_9_cnu_40_in_1, msg_to_check_it_9_cnu_40_in_2, msg_to_check_it_9_cnu_40_in_3, msg_to_check_it_9_cnu_40_in_4, msg_to_check_it_9_cnu_40_in_5, msg_to_check_it_9_cnu_41_in_0, msg_to_check_it_9_cnu_41_in_1, msg_to_check_it_9_cnu_41_in_2, msg_to_check_it_9_cnu_41_in_3, msg_to_check_it_9_cnu_41_in_4, msg_to_check_it_9_cnu_41_in_5, msg_to_check_it_9_cnu_42_in_0, msg_to_check_it_9_cnu_42_in_1, msg_to_check_it_9_cnu_42_in_2, msg_to_check_it_9_cnu_42_in_3, msg_to_check_it_9_cnu_42_in_4, msg_to_check_it_9_cnu_42_in_5, msg_to_check_it_9_cnu_43_in_0, msg_to_check_it_9_cnu_43_in_1, msg_to_check_it_9_cnu_43_in_2, msg_to_check_it_9_cnu_43_in_3, msg_to_check_it_9_cnu_43_in_4, msg_to_check_it_9_cnu_43_in_5, msg_to_check_it_9_cnu_44_in_0, msg_to_check_it_9_cnu_44_in_1, msg_to_check_it_9_cnu_44_in_2, msg_to_check_it_9_cnu_44_in_3, msg_to_check_it_9_cnu_44_in_4, msg_to_check_it_9_cnu_44_in_5, msg_to_check_it_9_cnu_45_in_0, msg_to_check_it_9_cnu_45_in_1, msg_to_check_it_9_cnu_45_in_2, msg_to_check_it_9_cnu_45_in_3, msg_to_check_it_9_cnu_45_in_4, msg_to_check_it_9_cnu_45_in_5, msg_to_check_it_9_cnu_46_in_0, msg_to_check_it_9_cnu_46_in_1, msg_to_check_it_9_cnu_46_in_2, msg_to_check_it_9_cnu_46_in_3, msg_to_check_it_9_cnu_46_in_4, msg_to_check_it_9_cnu_46_in_5, msg_to_check_it_9_cnu_47_in_0, msg_to_check_it_9_cnu_47_in_1, msg_to_check_it_9_cnu_47_in_2, msg_to_check_it_9_cnu_47_in_3, msg_to_check_it_9_cnu_47_in_4, msg_to_check_it_9_cnu_47_in_5, msg_to_check_it_9_cnu_48_in_0, msg_to_check_it_9_cnu_48_in_1, msg_to_check_it_9_cnu_48_in_2, msg_to_check_it_9_cnu_48_in_3, msg_to_check_it_9_cnu_48_in_4, msg_to_check_it_9_cnu_48_in_5, msg_to_check_it_9_cnu_49_in_0, msg_to_check_it_9_cnu_49_in_1, msg_to_check_it_9_cnu_49_in_2, msg_to_check_it_9_cnu_49_in_3, msg_to_check_it_9_cnu_49_in_4, msg_to_check_it_9_cnu_49_in_5, msg_to_check_it_9_cnu_50_in_0, msg_to_check_it_9_cnu_50_in_1, msg_to_check_it_9_cnu_50_in_2, msg_to_check_it_9_cnu_50_in_3, msg_to_check_it_9_cnu_50_in_4, msg_to_check_it_9_cnu_50_in_5, msg_to_check_it_9_cnu_51_in_0, msg_to_check_it_9_cnu_51_in_1, msg_to_check_it_9_cnu_51_in_2, msg_to_check_it_9_cnu_51_in_3, msg_to_check_it_9_cnu_51_in_4, msg_to_check_it_9_cnu_51_in_5, msg_to_check_it_9_cnu_52_in_0, msg_to_check_it_9_cnu_52_in_1, msg_to_check_it_9_cnu_52_in_2, msg_to_check_it_9_cnu_52_in_3, msg_to_check_it_9_cnu_52_in_4, msg_to_check_it_9_cnu_52_in_5, msg_to_check_it_9_cnu_53_in_0, msg_to_check_it_9_cnu_53_in_1, msg_to_check_it_9_cnu_53_in_2, msg_to_check_it_9_cnu_53_in_3, msg_to_check_it_9_cnu_53_in_4, msg_to_check_it_9_cnu_53_in_5, msg_to_check_it_9_cnu_54_in_0, msg_to_check_it_9_cnu_54_in_1, msg_to_check_it_9_cnu_54_in_2, msg_to_check_it_9_cnu_54_in_3, msg_to_check_it_9_cnu_54_in_4, msg_to_check_it_9_cnu_54_in_5, msg_to_check_it_9_cnu_55_in_0, msg_to_check_it_9_cnu_55_in_1, msg_to_check_it_9_cnu_55_in_2, msg_to_check_it_9_cnu_55_in_3, msg_to_check_it_9_cnu_55_in_4, msg_to_check_it_9_cnu_55_in_5, msg_to_check_it_9_cnu_56_in_0, msg_to_check_it_9_cnu_56_in_1, msg_to_check_it_9_cnu_56_in_2, msg_to_check_it_9_cnu_56_in_3, msg_to_check_it_9_cnu_56_in_4, msg_to_check_it_9_cnu_56_in_5, msg_to_check_it_9_cnu_57_in_0, msg_to_check_it_9_cnu_57_in_1, msg_to_check_it_9_cnu_57_in_2, msg_to_check_it_9_cnu_57_in_3, msg_to_check_it_9_cnu_57_in_4, msg_to_check_it_9_cnu_57_in_5, msg_to_check_it_9_cnu_58_in_0, msg_to_check_it_9_cnu_58_in_1, msg_to_check_it_9_cnu_58_in_2, msg_to_check_it_9_cnu_58_in_3, msg_to_check_it_9_cnu_58_in_4, msg_to_check_it_9_cnu_58_in_5, msg_to_check_it_9_cnu_59_in_0, msg_to_check_it_9_cnu_59_in_1, msg_to_check_it_9_cnu_59_in_2, msg_to_check_it_9_cnu_59_in_3, msg_to_check_it_9_cnu_59_in_4, msg_to_check_it_9_cnu_59_in_5, msg_to_check_it_9_cnu_60_in_0, msg_to_check_it_9_cnu_60_in_1, msg_to_check_it_9_cnu_60_in_2, msg_to_check_it_9_cnu_60_in_3, msg_to_check_it_9_cnu_60_in_4, msg_to_check_it_9_cnu_60_in_5, msg_to_check_it_9_cnu_61_in_0, msg_to_check_it_9_cnu_61_in_1, msg_to_check_it_9_cnu_61_in_2, msg_to_check_it_9_cnu_61_in_3, msg_to_check_it_9_cnu_61_in_4, msg_to_check_it_9_cnu_61_in_5, msg_to_check_it_9_cnu_62_in_0, msg_to_check_it_9_cnu_62_in_1, msg_to_check_it_9_cnu_62_in_2, msg_to_check_it_9_cnu_62_in_3, msg_to_check_it_9_cnu_62_in_4, msg_to_check_it_9_cnu_62_in_5, msg_to_check_it_9_cnu_63_in_0, msg_to_check_it_9_cnu_63_in_1, msg_to_check_it_9_cnu_63_in_2, msg_to_check_it_9_cnu_63_in_3, msg_to_check_it_9_cnu_63_in_4, msg_to_check_it_9_cnu_63_in_5, msg_to_check_it_9_cnu_64_in_0, msg_to_check_it_9_cnu_64_in_1, msg_to_check_it_9_cnu_64_in_2, msg_to_check_it_9_cnu_64_in_3, msg_to_check_it_9_cnu_64_in_4, msg_to_check_it_9_cnu_64_in_5, msg_to_check_it_9_cnu_65_in_0, msg_to_check_it_9_cnu_65_in_1, msg_to_check_it_9_cnu_65_in_2, msg_to_check_it_9_cnu_65_in_3, msg_to_check_it_9_cnu_65_in_4, msg_to_check_it_9_cnu_65_in_5, msg_to_check_it_9_cnu_66_in_0, msg_to_check_it_9_cnu_66_in_1, msg_to_check_it_9_cnu_66_in_2, msg_to_check_it_9_cnu_66_in_3, msg_to_check_it_9_cnu_66_in_4, msg_to_check_it_9_cnu_66_in_5, msg_to_check_it_9_cnu_67_in_0, msg_to_check_it_9_cnu_67_in_1, msg_to_check_it_9_cnu_67_in_2, msg_to_check_it_9_cnu_67_in_3, msg_to_check_it_9_cnu_67_in_4, msg_to_check_it_9_cnu_67_in_5, msg_to_check_it_9_cnu_68_in_0, msg_to_check_it_9_cnu_68_in_1, msg_to_check_it_9_cnu_68_in_2, msg_to_check_it_9_cnu_68_in_3, msg_to_check_it_9_cnu_68_in_4, msg_to_check_it_9_cnu_68_in_5, msg_to_check_it_9_cnu_69_in_0, msg_to_check_it_9_cnu_69_in_1, msg_to_check_it_9_cnu_69_in_2, msg_to_check_it_9_cnu_69_in_3, msg_to_check_it_9_cnu_69_in_4, msg_to_check_it_9_cnu_69_in_5, msg_to_check_it_9_cnu_70_in_0, msg_to_check_it_9_cnu_70_in_1, msg_to_check_it_9_cnu_70_in_2, msg_to_check_it_9_cnu_70_in_3, msg_to_check_it_9_cnu_70_in_4, msg_to_check_it_9_cnu_70_in_5, msg_to_check_it_9_cnu_71_in_0, msg_to_check_it_9_cnu_71_in_1, msg_to_check_it_9_cnu_71_in_2, msg_to_check_it_9_cnu_71_in_3, msg_to_check_it_9_cnu_71_in_4, msg_to_check_it_9_cnu_71_in_5, msg_to_check_it_9_cnu_72_in_0, msg_to_check_it_9_cnu_72_in_1, msg_to_check_it_9_cnu_72_in_2, msg_to_check_it_9_cnu_72_in_3, msg_to_check_it_9_cnu_72_in_4, msg_to_check_it_9_cnu_72_in_5, msg_to_check_it_9_cnu_73_in_0, msg_to_check_it_9_cnu_73_in_1, msg_to_check_it_9_cnu_73_in_2, msg_to_check_it_9_cnu_73_in_3, msg_to_check_it_9_cnu_73_in_4, msg_to_check_it_9_cnu_73_in_5, msg_to_check_it_9_cnu_74_in_0, msg_to_check_it_9_cnu_74_in_1, msg_to_check_it_9_cnu_74_in_2, msg_to_check_it_9_cnu_74_in_3, msg_to_check_it_9_cnu_74_in_4, msg_to_check_it_9_cnu_74_in_5, msg_to_check_it_9_cnu_75_in_0, msg_to_check_it_9_cnu_75_in_1, msg_to_check_it_9_cnu_75_in_2, msg_to_check_it_9_cnu_75_in_3, msg_to_check_it_9_cnu_75_in_4, msg_to_check_it_9_cnu_75_in_5, msg_to_check_it_9_cnu_76_in_0, msg_to_check_it_9_cnu_76_in_1, msg_to_check_it_9_cnu_76_in_2, msg_to_check_it_9_cnu_76_in_3, msg_to_check_it_9_cnu_76_in_4, msg_to_check_it_9_cnu_76_in_5, msg_to_check_it_9_cnu_77_in_0, msg_to_check_it_9_cnu_77_in_1, msg_to_check_it_9_cnu_77_in_2, msg_to_check_it_9_cnu_77_in_3, msg_to_check_it_9_cnu_77_in_4, msg_to_check_it_9_cnu_77_in_5, msg_to_check_it_9_cnu_78_in_0, msg_to_check_it_9_cnu_78_in_1, msg_to_check_it_9_cnu_78_in_2, msg_to_check_it_9_cnu_78_in_3, msg_to_check_it_9_cnu_78_in_4, msg_to_check_it_9_cnu_78_in_5, msg_to_check_it_9_cnu_79_in_0, msg_to_check_it_9_cnu_79_in_1, msg_to_check_it_9_cnu_79_in_2, msg_to_check_it_9_cnu_79_in_3, msg_to_check_it_9_cnu_79_in_4, msg_to_check_it_9_cnu_79_in_5, msg_to_check_it_9_cnu_80_in_0, msg_to_check_it_9_cnu_80_in_1, msg_to_check_it_9_cnu_80_in_2, msg_to_check_it_9_cnu_80_in_3, msg_to_check_it_9_cnu_80_in_4, msg_to_check_it_9_cnu_80_in_5, msg_to_check_it_9_cnu_81_in_0, msg_to_check_it_9_cnu_81_in_1, msg_to_check_it_9_cnu_81_in_2, msg_to_check_it_9_cnu_81_in_3, msg_to_check_it_9_cnu_81_in_4, msg_to_check_it_9_cnu_81_in_5, msg_to_check_it_9_cnu_82_in_0, msg_to_check_it_9_cnu_82_in_1, msg_to_check_it_9_cnu_82_in_2, msg_to_check_it_9_cnu_82_in_3, msg_to_check_it_9_cnu_82_in_4, msg_to_check_it_9_cnu_82_in_5, msg_to_check_it_9_cnu_83_in_0, msg_to_check_it_9_cnu_83_in_1, msg_to_check_it_9_cnu_83_in_2, msg_to_check_it_9_cnu_83_in_3, msg_to_check_it_9_cnu_83_in_4, msg_to_check_it_9_cnu_83_in_5, msg_to_check_it_9_cnu_84_in_0, msg_to_check_it_9_cnu_84_in_1, msg_to_check_it_9_cnu_84_in_2, msg_to_check_it_9_cnu_84_in_3, msg_to_check_it_9_cnu_84_in_4, msg_to_check_it_9_cnu_84_in_5, msg_to_check_it_9_cnu_85_in_0, msg_to_check_it_9_cnu_85_in_1, msg_to_check_it_9_cnu_85_in_2, msg_to_check_it_9_cnu_85_in_3, msg_to_check_it_9_cnu_85_in_4, msg_to_check_it_9_cnu_85_in_5, msg_to_check_it_9_cnu_86_in_0, msg_to_check_it_9_cnu_86_in_1, msg_to_check_it_9_cnu_86_in_2, msg_to_check_it_9_cnu_86_in_3, msg_to_check_it_9_cnu_86_in_4, msg_to_check_it_9_cnu_86_in_5, msg_to_check_it_9_cnu_87_in_0, msg_to_check_it_9_cnu_87_in_1, msg_to_check_it_9_cnu_87_in_2, msg_to_check_it_9_cnu_87_in_3, msg_to_check_it_9_cnu_87_in_4, msg_to_check_it_9_cnu_87_in_5, msg_to_check_it_9_cnu_88_in_0, msg_to_check_it_9_cnu_88_in_1, msg_to_check_it_9_cnu_88_in_2, msg_to_check_it_9_cnu_88_in_3, msg_to_check_it_9_cnu_88_in_4, msg_to_check_it_9_cnu_88_in_5, msg_to_check_it_9_cnu_89_in_0, msg_to_check_it_9_cnu_89_in_1, msg_to_check_it_9_cnu_89_in_2, msg_to_check_it_9_cnu_89_in_3, msg_to_check_it_9_cnu_89_in_4, msg_to_check_it_9_cnu_89_in_5, msg_to_check_it_9_cnu_90_in_0, msg_to_check_it_9_cnu_90_in_1, msg_to_check_it_9_cnu_90_in_2, msg_to_check_it_9_cnu_90_in_3, msg_to_check_it_9_cnu_90_in_4, msg_to_check_it_9_cnu_90_in_5, msg_to_check_it_9_cnu_91_in_0, msg_to_check_it_9_cnu_91_in_1, msg_to_check_it_9_cnu_91_in_2, msg_to_check_it_9_cnu_91_in_3, msg_to_check_it_9_cnu_91_in_4, msg_to_check_it_9_cnu_91_in_5, msg_to_check_it_9_cnu_92_in_0, msg_to_check_it_9_cnu_92_in_1, msg_to_check_it_9_cnu_92_in_2, msg_to_check_it_9_cnu_92_in_3, msg_to_check_it_9_cnu_92_in_4, msg_to_check_it_9_cnu_92_in_5, msg_to_check_it_9_cnu_93_in_0, msg_to_check_it_9_cnu_93_in_1, msg_to_check_it_9_cnu_93_in_2, msg_to_check_it_9_cnu_93_in_3, msg_to_check_it_9_cnu_93_in_4, msg_to_check_it_9_cnu_93_in_5, msg_to_check_it_9_cnu_94_in_0, msg_to_check_it_9_cnu_94_in_1, msg_to_check_it_9_cnu_94_in_2, msg_to_check_it_9_cnu_94_in_3, msg_to_check_it_9_cnu_94_in_4, msg_to_check_it_9_cnu_94_in_5, msg_to_check_it_9_cnu_95_in_0, msg_to_check_it_9_cnu_95_in_1, msg_to_check_it_9_cnu_95_in_2, msg_to_check_it_9_cnu_95_in_3, msg_to_check_it_9_cnu_95_in_4, msg_to_check_it_9_cnu_95_in_5, msg_to_check_it_9_cnu_96_in_0, msg_to_check_it_9_cnu_96_in_1, msg_to_check_it_9_cnu_96_in_2, msg_to_check_it_9_cnu_96_in_3, msg_to_check_it_9_cnu_96_in_4, msg_to_check_it_9_cnu_96_in_5, msg_to_check_it_9_cnu_97_in_0, msg_to_check_it_9_cnu_97_in_1, msg_to_check_it_9_cnu_97_in_2, msg_to_check_it_9_cnu_97_in_3, msg_to_check_it_9_cnu_97_in_4, msg_to_check_it_9_cnu_97_in_5, msg_to_check_it_9_cnu_98_in_0, msg_to_check_it_9_cnu_98_in_1, msg_to_check_it_9_cnu_98_in_2, msg_to_check_it_9_cnu_98_in_3, msg_to_check_it_9_cnu_98_in_4, msg_to_check_it_9_cnu_98_in_5, msg_to_check_it_10_cnu_0_in_0, msg_to_check_it_10_cnu_0_in_1, msg_to_check_it_10_cnu_0_in_2, msg_to_check_it_10_cnu_0_in_3, msg_to_check_it_10_cnu_0_in_4, msg_to_check_it_10_cnu_0_in_5, msg_to_check_it_10_cnu_1_in_0, msg_to_check_it_10_cnu_1_in_1, msg_to_check_it_10_cnu_1_in_2, msg_to_check_it_10_cnu_1_in_3, msg_to_check_it_10_cnu_1_in_4, msg_to_check_it_10_cnu_1_in_5, msg_to_check_it_10_cnu_2_in_0, msg_to_check_it_10_cnu_2_in_1, msg_to_check_it_10_cnu_2_in_2, msg_to_check_it_10_cnu_2_in_3, msg_to_check_it_10_cnu_2_in_4, msg_to_check_it_10_cnu_2_in_5, msg_to_check_it_10_cnu_3_in_0, msg_to_check_it_10_cnu_3_in_1, msg_to_check_it_10_cnu_3_in_2, msg_to_check_it_10_cnu_3_in_3, msg_to_check_it_10_cnu_3_in_4, msg_to_check_it_10_cnu_3_in_5, msg_to_check_it_10_cnu_4_in_0, msg_to_check_it_10_cnu_4_in_1, msg_to_check_it_10_cnu_4_in_2, msg_to_check_it_10_cnu_4_in_3, msg_to_check_it_10_cnu_4_in_4, msg_to_check_it_10_cnu_4_in_5, msg_to_check_it_10_cnu_5_in_0, msg_to_check_it_10_cnu_5_in_1, msg_to_check_it_10_cnu_5_in_2, msg_to_check_it_10_cnu_5_in_3, msg_to_check_it_10_cnu_5_in_4, msg_to_check_it_10_cnu_5_in_5, msg_to_check_it_10_cnu_6_in_0, msg_to_check_it_10_cnu_6_in_1, msg_to_check_it_10_cnu_6_in_2, msg_to_check_it_10_cnu_6_in_3, msg_to_check_it_10_cnu_6_in_4, msg_to_check_it_10_cnu_6_in_5, msg_to_check_it_10_cnu_7_in_0, msg_to_check_it_10_cnu_7_in_1, msg_to_check_it_10_cnu_7_in_2, msg_to_check_it_10_cnu_7_in_3, msg_to_check_it_10_cnu_7_in_4, msg_to_check_it_10_cnu_7_in_5, msg_to_check_it_10_cnu_8_in_0, msg_to_check_it_10_cnu_8_in_1, msg_to_check_it_10_cnu_8_in_2, msg_to_check_it_10_cnu_8_in_3, msg_to_check_it_10_cnu_8_in_4, msg_to_check_it_10_cnu_8_in_5, msg_to_check_it_10_cnu_9_in_0, msg_to_check_it_10_cnu_9_in_1, msg_to_check_it_10_cnu_9_in_2, msg_to_check_it_10_cnu_9_in_3, msg_to_check_it_10_cnu_9_in_4, msg_to_check_it_10_cnu_9_in_5, msg_to_check_it_10_cnu_10_in_0, msg_to_check_it_10_cnu_10_in_1, msg_to_check_it_10_cnu_10_in_2, msg_to_check_it_10_cnu_10_in_3, msg_to_check_it_10_cnu_10_in_4, msg_to_check_it_10_cnu_10_in_5, msg_to_check_it_10_cnu_11_in_0, msg_to_check_it_10_cnu_11_in_1, msg_to_check_it_10_cnu_11_in_2, msg_to_check_it_10_cnu_11_in_3, msg_to_check_it_10_cnu_11_in_4, msg_to_check_it_10_cnu_11_in_5, msg_to_check_it_10_cnu_12_in_0, msg_to_check_it_10_cnu_12_in_1, msg_to_check_it_10_cnu_12_in_2, msg_to_check_it_10_cnu_12_in_3, msg_to_check_it_10_cnu_12_in_4, msg_to_check_it_10_cnu_12_in_5, msg_to_check_it_10_cnu_13_in_0, msg_to_check_it_10_cnu_13_in_1, msg_to_check_it_10_cnu_13_in_2, msg_to_check_it_10_cnu_13_in_3, msg_to_check_it_10_cnu_13_in_4, msg_to_check_it_10_cnu_13_in_5, msg_to_check_it_10_cnu_14_in_0, msg_to_check_it_10_cnu_14_in_1, msg_to_check_it_10_cnu_14_in_2, msg_to_check_it_10_cnu_14_in_3, msg_to_check_it_10_cnu_14_in_4, msg_to_check_it_10_cnu_14_in_5, msg_to_check_it_10_cnu_15_in_0, msg_to_check_it_10_cnu_15_in_1, msg_to_check_it_10_cnu_15_in_2, msg_to_check_it_10_cnu_15_in_3, msg_to_check_it_10_cnu_15_in_4, msg_to_check_it_10_cnu_15_in_5, msg_to_check_it_10_cnu_16_in_0, msg_to_check_it_10_cnu_16_in_1, msg_to_check_it_10_cnu_16_in_2, msg_to_check_it_10_cnu_16_in_3, msg_to_check_it_10_cnu_16_in_4, msg_to_check_it_10_cnu_16_in_5, msg_to_check_it_10_cnu_17_in_0, msg_to_check_it_10_cnu_17_in_1, msg_to_check_it_10_cnu_17_in_2, msg_to_check_it_10_cnu_17_in_3, msg_to_check_it_10_cnu_17_in_4, msg_to_check_it_10_cnu_17_in_5, msg_to_check_it_10_cnu_18_in_0, msg_to_check_it_10_cnu_18_in_1, msg_to_check_it_10_cnu_18_in_2, msg_to_check_it_10_cnu_18_in_3, msg_to_check_it_10_cnu_18_in_4, msg_to_check_it_10_cnu_18_in_5, msg_to_check_it_10_cnu_19_in_0, msg_to_check_it_10_cnu_19_in_1, msg_to_check_it_10_cnu_19_in_2, msg_to_check_it_10_cnu_19_in_3, msg_to_check_it_10_cnu_19_in_4, msg_to_check_it_10_cnu_19_in_5, msg_to_check_it_10_cnu_20_in_0, msg_to_check_it_10_cnu_20_in_1, msg_to_check_it_10_cnu_20_in_2, msg_to_check_it_10_cnu_20_in_3, msg_to_check_it_10_cnu_20_in_4, msg_to_check_it_10_cnu_20_in_5, msg_to_check_it_10_cnu_21_in_0, msg_to_check_it_10_cnu_21_in_1, msg_to_check_it_10_cnu_21_in_2, msg_to_check_it_10_cnu_21_in_3, msg_to_check_it_10_cnu_21_in_4, msg_to_check_it_10_cnu_21_in_5, msg_to_check_it_10_cnu_22_in_0, msg_to_check_it_10_cnu_22_in_1, msg_to_check_it_10_cnu_22_in_2, msg_to_check_it_10_cnu_22_in_3, msg_to_check_it_10_cnu_22_in_4, msg_to_check_it_10_cnu_22_in_5, msg_to_check_it_10_cnu_23_in_0, msg_to_check_it_10_cnu_23_in_1, msg_to_check_it_10_cnu_23_in_2, msg_to_check_it_10_cnu_23_in_3, msg_to_check_it_10_cnu_23_in_4, msg_to_check_it_10_cnu_23_in_5, msg_to_check_it_10_cnu_24_in_0, msg_to_check_it_10_cnu_24_in_1, msg_to_check_it_10_cnu_24_in_2, msg_to_check_it_10_cnu_24_in_3, msg_to_check_it_10_cnu_24_in_4, msg_to_check_it_10_cnu_24_in_5, msg_to_check_it_10_cnu_25_in_0, msg_to_check_it_10_cnu_25_in_1, msg_to_check_it_10_cnu_25_in_2, msg_to_check_it_10_cnu_25_in_3, msg_to_check_it_10_cnu_25_in_4, msg_to_check_it_10_cnu_25_in_5, msg_to_check_it_10_cnu_26_in_0, msg_to_check_it_10_cnu_26_in_1, msg_to_check_it_10_cnu_26_in_2, msg_to_check_it_10_cnu_26_in_3, msg_to_check_it_10_cnu_26_in_4, msg_to_check_it_10_cnu_26_in_5, msg_to_check_it_10_cnu_27_in_0, msg_to_check_it_10_cnu_27_in_1, msg_to_check_it_10_cnu_27_in_2, msg_to_check_it_10_cnu_27_in_3, msg_to_check_it_10_cnu_27_in_4, msg_to_check_it_10_cnu_27_in_5, msg_to_check_it_10_cnu_28_in_0, msg_to_check_it_10_cnu_28_in_1, msg_to_check_it_10_cnu_28_in_2, msg_to_check_it_10_cnu_28_in_3, msg_to_check_it_10_cnu_28_in_4, msg_to_check_it_10_cnu_28_in_5, msg_to_check_it_10_cnu_29_in_0, msg_to_check_it_10_cnu_29_in_1, msg_to_check_it_10_cnu_29_in_2, msg_to_check_it_10_cnu_29_in_3, msg_to_check_it_10_cnu_29_in_4, msg_to_check_it_10_cnu_29_in_5, msg_to_check_it_10_cnu_30_in_0, msg_to_check_it_10_cnu_30_in_1, msg_to_check_it_10_cnu_30_in_2, msg_to_check_it_10_cnu_30_in_3, msg_to_check_it_10_cnu_30_in_4, msg_to_check_it_10_cnu_30_in_5, msg_to_check_it_10_cnu_31_in_0, msg_to_check_it_10_cnu_31_in_1, msg_to_check_it_10_cnu_31_in_2, msg_to_check_it_10_cnu_31_in_3, msg_to_check_it_10_cnu_31_in_4, msg_to_check_it_10_cnu_31_in_5, msg_to_check_it_10_cnu_32_in_0, msg_to_check_it_10_cnu_32_in_1, msg_to_check_it_10_cnu_32_in_2, msg_to_check_it_10_cnu_32_in_3, msg_to_check_it_10_cnu_32_in_4, msg_to_check_it_10_cnu_32_in_5, msg_to_check_it_10_cnu_33_in_0, msg_to_check_it_10_cnu_33_in_1, msg_to_check_it_10_cnu_33_in_2, msg_to_check_it_10_cnu_33_in_3, msg_to_check_it_10_cnu_33_in_4, msg_to_check_it_10_cnu_33_in_5, msg_to_check_it_10_cnu_34_in_0, msg_to_check_it_10_cnu_34_in_1, msg_to_check_it_10_cnu_34_in_2, msg_to_check_it_10_cnu_34_in_3, msg_to_check_it_10_cnu_34_in_4, msg_to_check_it_10_cnu_34_in_5, msg_to_check_it_10_cnu_35_in_0, msg_to_check_it_10_cnu_35_in_1, msg_to_check_it_10_cnu_35_in_2, msg_to_check_it_10_cnu_35_in_3, msg_to_check_it_10_cnu_35_in_4, msg_to_check_it_10_cnu_35_in_5, msg_to_check_it_10_cnu_36_in_0, msg_to_check_it_10_cnu_36_in_1, msg_to_check_it_10_cnu_36_in_2, msg_to_check_it_10_cnu_36_in_3, msg_to_check_it_10_cnu_36_in_4, msg_to_check_it_10_cnu_36_in_5, msg_to_check_it_10_cnu_37_in_0, msg_to_check_it_10_cnu_37_in_1, msg_to_check_it_10_cnu_37_in_2, msg_to_check_it_10_cnu_37_in_3, msg_to_check_it_10_cnu_37_in_4, msg_to_check_it_10_cnu_37_in_5, msg_to_check_it_10_cnu_38_in_0, msg_to_check_it_10_cnu_38_in_1, msg_to_check_it_10_cnu_38_in_2, msg_to_check_it_10_cnu_38_in_3, msg_to_check_it_10_cnu_38_in_4, msg_to_check_it_10_cnu_38_in_5, msg_to_check_it_10_cnu_39_in_0, msg_to_check_it_10_cnu_39_in_1, msg_to_check_it_10_cnu_39_in_2, msg_to_check_it_10_cnu_39_in_3, msg_to_check_it_10_cnu_39_in_4, msg_to_check_it_10_cnu_39_in_5, msg_to_check_it_10_cnu_40_in_0, msg_to_check_it_10_cnu_40_in_1, msg_to_check_it_10_cnu_40_in_2, msg_to_check_it_10_cnu_40_in_3, msg_to_check_it_10_cnu_40_in_4, msg_to_check_it_10_cnu_40_in_5, msg_to_check_it_10_cnu_41_in_0, msg_to_check_it_10_cnu_41_in_1, msg_to_check_it_10_cnu_41_in_2, msg_to_check_it_10_cnu_41_in_3, msg_to_check_it_10_cnu_41_in_4, msg_to_check_it_10_cnu_41_in_5, msg_to_check_it_10_cnu_42_in_0, msg_to_check_it_10_cnu_42_in_1, msg_to_check_it_10_cnu_42_in_2, msg_to_check_it_10_cnu_42_in_3, msg_to_check_it_10_cnu_42_in_4, msg_to_check_it_10_cnu_42_in_5, msg_to_check_it_10_cnu_43_in_0, msg_to_check_it_10_cnu_43_in_1, msg_to_check_it_10_cnu_43_in_2, msg_to_check_it_10_cnu_43_in_3, msg_to_check_it_10_cnu_43_in_4, msg_to_check_it_10_cnu_43_in_5, msg_to_check_it_10_cnu_44_in_0, msg_to_check_it_10_cnu_44_in_1, msg_to_check_it_10_cnu_44_in_2, msg_to_check_it_10_cnu_44_in_3, msg_to_check_it_10_cnu_44_in_4, msg_to_check_it_10_cnu_44_in_5, msg_to_check_it_10_cnu_45_in_0, msg_to_check_it_10_cnu_45_in_1, msg_to_check_it_10_cnu_45_in_2, msg_to_check_it_10_cnu_45_in_3, msg_to_check_it_10_cnu_45_in_4, msg_to_check_it_10_cnu_45_in_5, msg_to_check_it_10_cnu_46_in_0, msg_to_check_it_10_cnu_46_in_1, msg_to_check_it_10_cnu_46_in_2, msg_to_check_it_10_cnu_46_in_3, msg_to_check_it_10_cnu_46_in_4, msg_to_check_it_10_cnu_46_in_5, msg_to_check_it_10_cnu_47_in_0, msg_to_check_it_10_cnu_47_in_1, msg_to_check_it_10_cnu_47_in_2, msg_to_check_it_10_cnu_47_in_3, msg_to_check_it_10_cnu_47_in_4, msg_to_check_it_10_cnu_47_in_5, msg_to_check_it_10_cnu_48_in_0, msg_to_check_it_10_cnu_48_in_1, msg_to_check_it_10_cnu_48_in_2, msg_to_check_it_10_cnu_48_in_3, msg_to_check_it_10_cnu_48_in_4, msg_to_check_it_10_cnu_48_in_5, msg_to_check_it_10_cnu_49_in_0, msg_to_check_it_10_cnu_49_in_1, msg_to_check_it_10_cnu_49_in_2, msg_to_check_it_10_cnu_49_in_3, msg_to_check_it_10_cnu_49_in_4, msg_to_check_it_10_cnu_49_in_5, msg_to_check_it_10_cnu_50_in_0, msg_to_check_it_10_cnu_50_in_1, msg_to_check_it_10_cnu_50_in_2, msg_to_check_it_10_cnu_50_in_3, msg_to_check_it_10_cnu_50_in_4, msg_to_check_it_10_cnu_50_in_5, msg_to_check_it_10_cnu_51_in_0, msg_to_check_it_10_cnu_51_in_1, msg_to_check_it_10_cnu_51_in_2, msg_to_check_it_10_cnu_51_in_3, msg_to_check_it_10_cnu_51_in_4, msg_to_check_it_10_cnu_51_in_5, msg_to_check_it_10_cnu_52_in_0, msg_to_check_it_10_cnu_52_in_1, msg_to_check_it_10_cnu_52_in_2, msg_to_check_it_10_cnu_52_in_3, msg_to_check_it_10_cnu_52_in_4, msg_to_check_it_10_cnu_52_in_5, msg_to_check_it_10_cnu_53_in_0, msg_to_check_it_10_cnu_53_in_1, msg_to_check_it_10_cnu_53_in_2, msg_to_check_it_10_cnu_53_in_3, msg_to_check_it_10_cnu_53_in_4, msg_to_check_it_10_cnu_53_in_5, msg_to_check_it_10_cnu_54_in_0, msg_to_check_it_10_cnu_54_in_1, msg_to_check_it_10_cnu_54_in_2, msg_to_check_it_10_cnu_54_in_3, msg_to_check_it_10_cnu_54_in_4, msg_to_check_it_10_cnu_54_in_5, msg_to_check_it_10_cnu_55_in_0, msg_to_check_it_10_cnu_55_in_1, msg_to_check_it_10_cnu_55_in_2, msg_to_check_it_10_cnu_55_in_3, msg_to_check_it_10_cnu_55_in_4, msg_to_check_it_10_cnu_55_in_5, msg_to_check_it_10_cnu_56_in_0, msg_to_check_it_10_cnu_56_in_1, msg_to_check_it_10_cnu_56_in_2, msg_to_check_it_10_cnu_56_in_3, msg_to_check_it_10_cnu_56_in_4, msg_to_check_it_10_cnu_56_in_5, msg_to_check_it_10_cnu_57_in_0, msg_to_check_it_10_cnu_57_in_1, msg_to_check_it_10_cnu_57_in_2, msg_to_check_it_10_cnu_57_in_3, msg_to_check_it_10_cnu_57_in_4, msg_to_check_it_10_cnu_57_in_5, msg_to_check_it_10_cnu_58_in_0, msg_to_check_it_10_cnu_58_in_1, msg_to_check_it_10_cnu_58_in_2, msg_to_check_it_10_cnu_58_in_3, msg_to_check_it_10_cnu_58_in_4, msg_to_check_it_10_cnu_58_in_5, msg_to_check_it_10_cnu_59_in_0, msg_to_check_it_10_cnu_59_in_1, msg_to_check_it_10_cnu_59_in_2, msg_to_check_it_10_cnu_59_in_3, msg_to_check_it_10_cnu_59_in_4, msg_to_check_it_10_cnu_59_in_5, msg_to_check_it_10_cnu_60_in_0, msg_to_check_it_10_cnu_60_in_1, msg_to_check_it_10_cnu_60_in_2, msg_to_check_it_10_cnu_60_in_3, msg_to_check_it_10_cnu_60_in_4, msg_to_check_it_10_cnu_60_in_5, msg_to_check_it_10_cnu_61_in_0, msg_to_check_it_10_cnu_61_in_1, msg_to_check_it_10_cnu_61_in_2, msg_to_check_it_10_cnu_61_in_3, msg_to_check_it_10_cnu_61_in_4, msg_to_check_it_10_cnu_61_in_5, msg_to_check_it_10_cnu_62_in_0, msg_to_check_it_10_cnu_62_in_1, msg_to_check_it_10_cnu_62_in_2, msg_to_check_it_10_cnu_62_in_3, msg_to_check_it_10_cnu_62_in_4, msg_to_check_it_10_cnu_62_in_5, msg_to_check_it_10_cnu_63_in_0, msg_to_check_it_10_cnu_63_in_1, msg_to_check_it_10_cnu_63_in_2, msg_to_check_it_10_cnu_63_in_3, msg_to_check_it_10_cnu_63_in_4, msg_to_check_it_10_cnu_63_in_5, msg_to_check_it_10_cnu_64_in_0, msg_to_check_it_10_cnu_64_in_1, msg_to_check_it_10_cnu_64_in_2, msg_to_check_it_10_cnu_64_in_3, msg_to_check_it_10_cnu_64_in_4, msg_to_check_it_10_cnu_64_in_5, msg_to_check_it_10_cnu_65_in_0, msg_to_check_it_10_cnu_65_in_1, msg_to_check_it_10_cnu_65_in_2, msg_to_check_it_10_cnu_65_in_3, msg_to_check_it_10_cnu_65_in_4, msg_to_check_it_10_cnu_65_in_5, msg_to_check_it_10_cnu_66_in_0, msg_to_check_it_10_cnu_66_in_1, msg_to_check_it_10_cnu_66_in_2, msg_to_check_it_10_cnu_66_in_3, msg_to_check_it_10_cnu_66_in_4, msg_to_check_it_10_cnu_66_in_5, msg_to_check_it_10_cnu_67_in_0, msg_to_check_it_10_cnu_67_in_1, msg_to_check_it_10_cnu_67_in_2, msg_to_check_it_10_cnu_67_in_3, msg_to_check_it_10_cnu_67_in_4, msg_to_check_it_10_cnu_67_in_5, msg_to_check_it_10_cnu_68_in_0, msg_to_check_it_10_cnu_68_in_1, msg_to_check_it_10_cnu_68_in_2, msg_to_check_it_10_cnu_68_in_3, msg_to_check_it_10_cnu_68_in_4, msg_to_check_it_10_cnu_68_in_5, msg_to_check_it_10_cnu_69_in_0, msg_to_check_it_10_cnu_69_in_1, msg_to_check_it_10_cnu_69_in_2, msg_to_check_it_10_cnu_69_in_3, msg_to_check_it_10_cnu_69_in_4, msg_to_check_it_10_cnu_69_in_5, msg_to_check_it_10_cnu_70_in_0, msg_to_check_it_10_cnu_70_in_1, msg_to_check_it_10_cnu_70_in_2, msg_to_check_it_10_cnu_70_in_3, msg_to_check_it_10_cnu_70_in_4, msg_to_check_it_10_cnu_70_in_5, msg_to_check_it_10_cnu_71_in_0, msg_to_check_it_10_cnu_71_in_1, msg_to_check_it_10_cnu_71_in_2, msg_to_check_it_10_cnu_71_in_3, msg_to_check_it_10_cnu_71_in_4, msg_to_check_it_10_cnu_71_in_5, msg_to_check_it_10_cnu_72_in_0, msg_to_check_it_10_cnu_72_in_1, msg_to_check_it_10_cnu_72_in_2, msg_to_check_it_10_cnu_72_in_3, msg_to_check_it_10_cnu_72_in_4, msg_to_check_it_10_cnu_72_in_5, msg_to_check_it_10_cnu_73_in_0, msg_to_check_it_10_cnu_73_in_1, msg_to_check_it_10_cnu_73_in_2, msg_to_check_it_10_cnu_73_in_3, msg_to_check_it_10_cnu_73_in_4, msg_to_check_it_10_cnu_73_in_5, msg_to_check_it_10_cnu_74_in_0, msg_to_check_it_10_cnu_74_in_1, msg_to_check_it_10_cnu_74_in_2, msg_to_check_it_10_cnu_74_in_3, msg_to_check_it_10_cnu_74_in_4, msg_to_check_it_10_cnu_74_in_5, msg_to_check_it_10_cnu_75_in_0, msg_to_check_it_10_cnu_75_in_1, msg_to_check_it_10_cnu_75_in_2, msg_to_check_it_10_cnu_75_in_3, msg_to_check_it_10_cnu_75_in_4, msg_to_check_it_10_cnu_75_in_5, msg_to_check_it_10_cnu_76_in_0, msg_to_check_it_10_cnu_76_in_1, msg_to_check_it_10_cnu_76_in_2, msg_to_check_it_10_cnu_76_in_3, msg_to_check_it_10_cnu_76_in_4, msg_to_check_it_10_cnu_76_in_5, msg_to_check_it_10_cnu_77_in_0, msg_to_check_it_10_cnu_77_in_1, msg_to_check_it_10_cnu_77_in_2, msg_to_check_it_10_cnu_77_in_3, msg_to_check_it_10_cnu_77_in_4, msg_to_check_it_10_cnu_77_in_5, msg_to_check_it_10_cnu_78_in_0, msg_to_check_it_10_cnu_78_in_1, msg_to_check_it_10_cnu_78_in_2, msg_to_check_it_10_cnu_78_in_3, msg_to_check_it_10_cnu_78_in_4, msg_to_check_it_10_cnu_78_in_5, msg_to_check_it_10_cnu_79_in_0, msg_to_check_it_10_cnu_79_in_1, msg_to_check_it_10_cnu_79_in_2, msg_to_check_it_10_cnu_79_in_3, msg_to_check_it_10_cnu_79_in_4, msg_to_check_it_10_cnu_79_in_5, msg_to_check_it_10_cnu_80_in_0, msg_to_check_it_10_cnu_80_in_1, msg_to_check_it_10_cnu_80_in_2, msg_to_check_it_10_cnu_80_in_3, msg_to_check_it_10_cnu_80_in_4, msg_to_check_it_10_cnu_80_in_5, msg_to_check_it_10_cnu_81_in_0, msg_to_check_it_10_cnu_81_in_1, msg_to_check_it_10_cnu_81_in_2, msg_to_check_it_10_cnu_81_in_3, msg_to_check_it_10_cnu_81_in_4, msg_to_check_it_10_cnu_81_in_5, msg_to_check_it_10_cnu_82_in_0, msg_to_check_it_10_cnu_82_in_1, msg_to_check_it_10_cnu_82_in_2, msg_to_check_it_10_cnu_82_in_3, msg_to_check_it_10_cnu_82_in_4, msg_to_check_it_10_cnu_82_in_5, msg_to_check_it_10_cnu_83_in_0, msg_to_check_it_10_cnu_83_in_1, msg_to_check_it_10_cnu_83_in_2, msg_to_check_it_10_cnu_83_in_3, msg_to_check_it_10_cnu_83_in_4, msg_to_check_it_10_cnu_83_in_5, msg_to_check_it_10_cnu_84_in_0, msg_to_check_it_10_cnu_84_in_1, msg_to_check_it_10_cnu_84_in_2, msg_to_check_it_10_cnu_84_in_3, msg_to_check_it_10_cnu_84_in_4, msg_to_check_it_10_cnu_84_in_5, msg_to_check_it_10_cnu_85_in_0, msg_to_check_it_10_cnu_85_in_1, msg_to_check_it_10_cnu_85_in_2, msg_to_check_it_10_cnu_85_in_3, msg_to_check_it_10_cnu_85_in_4, msg_to_check_it_10_cnu_85_in_5, msg_to_check_it_10_cnu_86_in_0, msg_to_check_it_10_cnu_86_in_1, msg_to_check_it_10_cnu_86_in_2, msg_to_check_it_10_cnu_86_in_3, msg_to_check_it_10_cnu_86_in_4, msg_to_check_it_10_cnu_86_in_5, msg_to_check_it_10_cnu_87_in_0, msg_to_check_it_10_cnu_87_in_1, msg_to_check_it_10_cnu_87_in_2, msg_to_check_it_10_cnu_87_in_3, msg_to_check_it_10_cnu_87_in_4, msg_to_check_it_10_cnu_87_in_5, msg_to_check_it_10_cnu_88_in_0, msg_to_check_it_10_cnu_88_in_1, msg_to_check_it_10_cnu_88_in_2, msg_to_check_it_10_cnu_88_in_3, msg_to_check_it_10_cnu_88_in_4, msg_to_check_it_10_cnu_88_in_5, msg_to_check_it_10_cnu_89_in_0, msg_to_check_it_10_cnu_89_in_1, msg_to_check_it_10_cnu_89_in_2, msg_to_check_it_10_cnu_89_in_3, msg_to_check_it_10_cnu_89_in_4, msg_to_check_it_10_cnu_89_in_5, msg_to_check_it_10_cnu_90_in_0, msg_to_check_it_10_cnu_90_in_1, msg_to_check_it_10_cnu_90_in_2, msg_to_check_it_10_cnu_90_in_3, msg_to_check_it_10_cnu_90_in_4, msg_to_check_it_10_cnu_90_in_5, msg_to_check_it_10_cnu_91_in_0, msg_to_check_it_10_cnu_91_in_1, msg_to_check_it_10_cnu_91_in_2, msg_to_check_it_10_cnu_91_in_3, msg_to_check_it_10_cnu_91_in_4, msg_to_check_it_10_cnu_91_in_5, msg_to_check_it_10_cnu_92_in_0, msg_to_check_it_10_cnu_92_in_1, msg_to_check_it_10_cnu_92_in_2, msg_to_check_it_10_cnu_92_in_3, msg_to_check_it_10_cnu_92_in_4, msg_to_check_it_10_cnu_92_in_5, msg_to_check_it_10_cnu_93_in_0, msg_to_check_it_10_cnu_93_in_1, msg_to_check_it_10_cnu_93_in_2, msg_to_check_it_10_cnu_93_in_3, msg_to_check_it_10_cnu_93_in_4, msg_to_check_it_10_cnu_93_in_5, msg_to_check_it_10_cnu_94_in_0, msg_to_check_it_10_cnu_94_in_1, msg_to_check_it_10_cnu_94_in_2, msg_to_check_it_10_cnu_94_in_3, msg_to_check_it_10_cnu_94_in_4, msg_to_check_it_10_cnu_94_in_5, msg_to_check_it_10_cnu_95_in_0, msg_to_check_it_10_cnu_95_in_1, msg_to_check_it_10_cnu_95_in_2, msg_to_check_it_10_cnu_95_in_3, msg_to_check_it_10_cnu_95_in_4, msg_to_check_it_10_cnu_95_in_5, msg_to_check_it_10_cnu_96_in_0, msg_to_check_it_10_cnu_96_in_1, msg_to_check_it_10_cnu_96_in_2, msg_to_check_it_10_cnu_96_in_3, msg_to_check_it_10_cnu_96_in_4, msg_to_check_it_10_cnu_96_in_5, msg_to_check_it_10_cnu_97_in_0, msg_to_check_it_10_cnu_97_in_1, msg_to_check_it_10_cnu_97_in_2, msg_to_check_it_10_cnu_97_in_3, msg_to_check_it_10_cnu_97_in_4, msg_to_check_it_10_cnu_97_in_5, msg_to_check_it_10_cnu_98_in_0, msg_to_check_it_10_cnu_98_in_1, msg_to_check_it_10_cnu_98_in_2, msg_to_check_it_10_cnu_98_in_3, msg_to_check_it_10_cnu_98_in_4, msg_to_check_it_10_cnu_98_in_5, msg_to_check_it_11_cnu_0_in_0, msg_to_check_it_11_cnu_0_in_1, msg_to_check_it_11_cnu_0_in_2, msg_to_check_it_11_cnu_0_in_3, msg_to_check_it_11_cnu_0_in_4, msg_to_check_it_11_cnu_0_in_5, msg_to_check_it_11_cnu_1_in_0, msg_to_check_it_11_cnu_1_in_1, msg_to_check_it_11_cnu_1_in_2, msg_to_check_it_11_cnu_1_in_3, msg_to_check_it_11_cnu_1_in_4, msg_to_check_it_11_cnu_1_in_5, msg_to_check_it_11_cnu_2_in_0, msg_to_check_it_11_cnu_2_in_1, msg_to_check_it_11_cnu_2_in_2, msg_to_check_it_11_cnu_2_in_3, msg_to_check_it_11_cnu_2_in_4, msg_to_check_it_11_cnu_2_in_5, msg_to_check_it_11_cnu_3_in_0, msg_to_check_it_11_cnu_3_in_1, msg_to_check_it_11_cnu_3_in_2, msg_to_check_it_11_cnu_3_in_3, msg_to_check_it_11_cnu_3_in_4, msg_to_check_it_11_cnu_3_in_5, msg_to_check_it_11_cnu_4_in_0, msg_to_check_it_11_cnu_4_in_1, msg_to_check_it_11_cnu_4_in_2, msg_to_check_it_11_cnu_4_in_3, msg_to_check_it_11_cnu_4_in_4, msg_to_check_it_11_cnu_4_in_5, msg_to_check_it_11_cnu_5_in_0, msg_to_check_it_11_cnu_5_in_1, msg_to_check_it_11_cnu_5_in_2, msg_to_check_it_11_cnu_5_in_3, msg_to_check_it_11_cnu_5_in_4, msg_to_check_it_11_cnu_5_in_5, msg_to_check_it_11_cnu_6_in_0, msg_to_check_it_11_cnu_6_in_1, msg_to_check_it_11_cnu_6_in_2, msg_to_check_it_11_cnu_6_in_3, msg_to_check_it_11_cnu_6_in_4, msg_to_check_it_11_cnu_6_in_5, msg_to_check_it_11_cnu_7_in_0, msg_to_check_it_11_cnu_7_in_1, msg_to_check_it_11_cnu_7_in_2, msg_to_check_it_11_cnu_7_in_3, msg_to_check_it_11_cnu_7_in_4, msg_to_check_it_11_cnu_7_in_5, msg_to_check_it_11_cnu_8_in_0, msg_to_check_it_11_cnu_8_in_1, msg_to_check_it_11_cnu_8_in_2, msg_to_check_it_11_cnu_8_in_3, msg_to_check_it_11_cnu_8_in_4, msg_to_check_it_11_cnu_8_in_5, msg_to_check_it_11_cnu_9_in_0, msg_to_check_it_11_cnu_9_in_1, msg_to_check_it_11_cnu_9_in_2, msg_to_check_it_11_cnu_9_in_3, msg_to_check_it_11_cnu_9_in_4, msg_to_check_it_11_cnu_9_in_5, msg_to_check_it_11_cnu_10_in_0, msg_to_check_it_11_cnu_10_in_1, msg_to_check_it_11_cnu_10_in_2, msg_to_check_it_11_cnu_10_in_3, msg_to_check_it_11_cnu_10_in_4, msg_to_check_it_11_cnu_10_in_5, msg_to_check_it_11_cnu_11_in_0, msg_to_check_it_11_cnu_11_in_1, msg_to_check_it_11_cnu_11_in_2, msg_to_check_it_11_cnu_11_in_3, msg_to_check_it_11_cnu_11_in_4, msg_to_check_it_11_cnu_11_in_5, msg_to_check_it_11_cnu_12_in_0, msg_to_check_it_11_cnu_12_in_1, msg_to_check_it_11_cnu_12_in_2, msg_to_check_it_11_cnu_12_in_3, msg_to_check_it_11_cnu_12_in_4, msg_to_check_it_11_cnu_12_in_5, msg_to_check_it_11_cnu_13_in_0, msg_to_check_it_11_cnu_13_in_1, msg_to_check_it_11_cnu_13_in_2, msg_to_check_it_11_cnu_13_in_3, msg_to_check_it_11_cnu_13_in_4, msg_to_check_it_11_cnu_13_in_5, msg_to_check_it_11_cnu_14_in_0, msg_to_check_it_11_cnu_14_in_1, msg_to_check_it_11_cnu_14_in_2, msg_to_check_it_11_cnu_14_in_3, msg_to_check_it_11_cnu_14_in_4, msg_to_check_it_11_cnu_14_in_5, msg_to_check_it_11_cnu_15_in_0, msg_to_check_it_11_cnu_15_in_1, msg_to_check_it_11_cnu_15_in_2, msg_to_check_it_11_cnu_15_in_3, msg_to_check_it_11_cnu_15_in_4, msg_to_check_it_11_cnu_15_in_5, msg_to_check_it_11_cnu_16_in_0, msg_to_check_it_11_cnu_16_in_1, msg_to_check_it_11_cnu_16_in_2, msg_to_check_it_11_cnu_16_in_3, msg_to_check_it_11_cnu_16_in_4, msg_to_check_it_11_cnu_16_in_5, msg_to_check_it_11_cnu_17_in_0, msg_to_check_it_11_cnu_17_in_1, msg_to_check_it_11_cnu_17_in_2, msg_to_check_it_11_cnu_17_in_3, msg_to_check_it_11_cnu_17_in_4, msg_to_check_it_11_cnu_17_in_5, msg_to_check_it_11_cnu_18_in_0, msg_to_check_it_11_cnu_18_in_1, msg_to_check_it_11_cnu_18_in_2, msg_to_check_it_11_cnu_18_in_3, msg_to_check_it_11_cnu_18_in_4, msg_to_check_it_11_cnu_18_in_5, msg_to_check_it_11_cnu_19_in_0, msg_to_check_it_11_cnu_19_in_1, msg_to_check_it_11_cnu_19_in_2, msg_to_check_it_11_cnu_19_in_3, msg_to_check_it_11_cnu_19_in_4, msg_to_check_it_11_cnu_19_in_5, msg_to_check_it_11_cnu_20_in_0, msg_to_check_it_11_cnu_20_in_1, msg_to_check_it_11_cnu_20_in_2, msg_to_check_it_11_cnu_20_in_3, msg_to_check_it_11_cnu_20_in_4, msg_to_check_it_11_cnu_20_in_5, msg_to_check_it_11_cnu_21_in_0, msg_to_check_it_11_cnu_21_in_1, msg_to_check_it_11_cnu_21_in_2, msg_to_check_it_11_cnu_21_in_3, msg_to_check_it_11_cnu_21_in_4, msg_to_check_it_11_cnu_21_in_5, msg_to_check_it_11_cnu_22_in_0, msg_to_check_it_11_cnu_22_in_1, msg_to_check_it_11_cnu_22_in_2, msg_to_check_it_11_cnu_22_in_3, msg_to_check_it_11_cnu_22_in_4, msg_to_check_it_11_cnu_22_in_5, msg_to_check_it_11_cnu_23_in_0, msg_to_check_it_11_cnu_23_in_1, msg_to_check_it_11_cnu_23_in_2, msg_to_check_it_11_cnu_23_in_3, msg_to_check_it_11_cnu_23_in_4, msg_to_check_it_11_cnu_23_in_5, msg_to_check_it_11_cnu_24_in_0, msg_to_check_it_11_cnu_24_in_1, msg_to_check_it_11_cnu_24_in_2, msg_to_check_it_11_cnu_24_in_3, msg_to_check_it_11_cnu_24_in_4, msg_to_check_it_11_cnu_24_in_5, msg_to_check_it_11_cnu_25_in_0, msg_to_check_it_11_cnu_25_in_1, msg_to_check_it_11_cnu_25_in_2, msg_to_check_it_11_cnu_25_in_3, msg_to_check_it_11_cnu_25_in_4, msg_to_check_it_11_cnu_25_in_5, msg_to_check_it_11_cnu_26_in_0, msg_to_check_it_11_cnu_26_in_1, msg_to_check_it_11_cnu_26_in_2, msg_to_check_it_11_cnu_26_in_3, msg_to_check_it_11_cnu_26_in_4, msg_to_check_it_11_cnu_26_in_5, msg_to_check_it_11_cnu_27_in_0, msg_to_check_it_11_cnu_27_in_1, msg_to_check_it_11_cnu_27_in_2, msg_to_check_it_11_cnu_27_in_3, msg_to_check_it_11_cnu_27_in_4, msg_to_check_it_11_cnu_27_in_5, msg_to_check_it_11_cnu_28_in_0, msg_to_check_it_11_cnu_28_in_1, msg_to_check_it_11_cnu_28_in_2, msg_to_check_it_11_cnu_28_in_3, msg_to_check_it_11_cnu_28_in_4, msg_to_check_it_11_cnu_28_in_5, msg_to_check_it_11_cnu_29_in_0, msg_to_check_it_11_cnu_29_in_1, msg_to_check_it_11_cnu_29_in_2, msg_to_check_it_11_cnu_29_in_3, msg_to_check_it_11_cnu_29_in_4, msg_to_check_it_11_cnu_29_in_5, msg_to_check_it_11_cnu_30_in_0, msg_to_check_it_11_cnu_30_in_1, msg_to_check_it_11_cnu_30_in_2, msg_to_check_it_11_cnu_30_in_3, msg_to_check_it_11_cnu_30_in_4, msg_to_check_it_11_cnu_30_in_5, msg_to_check_it_11_cnu_31_in_0, msg_to_check_it_11_cnu_31_in_1, msg_to_check_it_11_cnu_31_in_2, msg_to_check_it_11_cnu_31_in_3, msg_to_check_it_11_cnu_31_in_4, msg_to_check_it_11_cnu_31_in_5, msg_to_check_it_11_cnu_32_in_0, msg_to_check_it_11_cnu_32_in_1, msg_to_check_it_11_cnu_32_in_2, msg_to_check_it_11_cnu_32_in_3, msg_to_check_it_11_cnu_32_in_4, msg_to_check_it_11_cnu_32_in_5, msg_to_check_it_11_cnu_33_in_0, msg_to_check_it_11_cnu_33_in_1, msg_to_check_it_11_cnu_33_in_2, msg_to_check_it_11_cnu_33_in_3, msg_to_check_it_11_cnu_33_in_4, msg_to_check_it_11_cnu_33_in_5, msg_to_check_it_11_cnu_34_in_0, msg_to_check_it_11_cnu_34_in_1, msg_to_check_it_11_cnu_34_in_2, msg_to_check_it_11_cnu_34_in_3, msg_to_check_it_11_cnu_34_in_4, msg_to_check_it_11_cnu_34_in_5, msg_to_check_it_11_cnu_35_in_0, msg_to_check_it_11_cnu_35_in_1, msg_to_check_it_11_cnu_35_in_2, msg_to_check_it_11_cnu_35_in_3, msg_to_check_it_11_cnu_35_in_4, msg_to_check_it_11_cnu_35_in_5, msg_to_check_it_11_cnu_36_in_0, msg_to_check_it_11_cnu_36_in_1, msg_to_check_it_11_cnu_36_in_2, msg_to_check_it_11_cnu_36_in_3, msg_to_check_it_11_cnu_36_in_4, msg_to_check_it_11_cnu_36_in_5, msg_to_check_it_11_cnu_37_in_0, msg_to_check_it_11_cnu_37_in_1, msg_to_check_it_11_cnu_37_in_2, msg_to_check_it_11_cnu_37_in_3, msg_to_check_it_11_cnu_37_in_4, msg_to_check_it_11_cnu_37_in_5, msg_to_check_it_11_cnu_38_in_0, msg_to_check_it_11_cnu_38_in_1, msg_to_check_it_11_cnu_38_in_2, msg_to_check_it_11_cnu_38_in_3, msg_to_check_it_11_cnu_38_in_4, msg_to_check_it_11_cnu_38_in_5, msg_to_check_it_11_cnu_39_in_0, msg_to_check_it_11_cnu_39_in_1, msg_to_check_it_11_cnu_39_in_2, msg_to_check_it_11_cnu_39_in_3, msg_to_check_it_11_cnu_39_in_4, msg_to_check_it_11_cnu_39_in_5, msg_to_check_it_11_cnu_40_in_0, msg_to_check_it_11_cnu_40_in_1, msg_to_check_it_11_cnu_40_in_2, msg_to_check_it_11_cnu_40_in_3, msg_to_check_it_11_cnu_40_in_4, msg_to_check_it_11_cnu_40_in_5, msg_to_check_it_11_cnu_41_in_0, msg_to_check_it_11_cnu_41_in_1, msg_to_check_it_11_cnu_41_in_2, msg_to_check_it_11_cnu_41_in_3, msg_to_check_it_11_cnu_41_in_4, msg_to_check_it_11_cnu_41_in_5, msg_to_check_it_11_cnu_42_in_0, msg_to_check_it_11_cnu_42_in_1, msg_to_check_it_11_cnu_42_in_2, msg_to_check_it_11_cnu_42_in_3, msg_to_check_it_11_cnu_42_in_4, msg_to_check_it_11_cnu_42_in_5, msg_to_check_it_11_cnu_43_in_0, msg_to_check_it_11_cnu_43_in_1, msg_to_check_it_11_cnu_43_in_2, msg_to_check_it_11_cnu_43_in_3, msg_to_check_it_11_cnu_43_in_4, msg_to_check_it_11_cnu_43_in_5, msg_to_check_it_11_cnu_44_in_0, msg_to_check_it_11_cnu_44_in_1, msg_to_check_it_11_cnu_44_in_2, msg_to_check_it_11_cnu_44_in_3, msg_to_check_it_11_cnu_44_in_4, msg_to_check_it_11_cnu_44_in_5, msg_to_check_it_11_cnu_45_in_0, msg_to_check_it_11_cnu_45_in_1, msg_to_check_it_11_cnu_45_in_2, msg_to_check_it_11_cnu_45_in_3, msg_to_check_it_11_cnu_45_in_4, msg_to_check_it_11_cnu_45_in_5, msg_to_check_it_11_cnu_46_in_0, msg_to_check_it_11_cnu_46_in_1, msg_to_check_it_11_cnu_46_in_2, msg_to_check_it_11_cnu_46_in_3, msg_to_check_it_11_cnu_46_in_4, msg_to_check_it_11_cnu_46_in_5, msg_to_check_it_11_cnu_47_in_0, msg_to_check_it_11_cnu_47_in_1, msg_to_check_it_11_cnu_47_in_2, msg_to_check_it_11_cnu_47_in_3, msg_to_check_it_11_cnu_47_in_4, msg_to_check_it_11_cnu_47_in_5, msg_to_check_it_11_cnu_48_in_0, msg_to_check_it_11_cnu_48_in_1, msg_to_check_it_11_cnu_48_in_2, msg_to_check_it_11_cnu_48_in_3, msg_to_check_it_11_cnu_48_in_4, msg_to_check_it_11_cnu_48_in_5, msg_to_check_it_11_cnu_49_in_0, msg_to_check_it_11_cnu_49_in_1, msg_to_check_it_11_cnu_49_in_2, msg_to_check_it_11_cnu_49_in_3, msg_to_check_it_11_cnu_49_in_4, msg_to_check_it_11_cnu_49_in_5, msg_to_check_it_11_cnu_50_in_0, msg_to_check_it_11_cnu_50_in_1, msg_to_check_it_11_cnu_50_in_2, msg_to_check_it_11_cnu_50_in_3, msg_to_check_it_11_cnu_50_in_4, msg_to_check_it_11_cnu_50_in_5, msg_to_check_it_11_cnu_51_in_0, msg_to_check_it_11_cnu_51_in_1, msg_to_check_it_11_cnu_51_in_2, msg_to_check_it_11_cnu_51_in_3, msg_to_check_it_11_cnu_51_in_4, msg_to_check_it_11_cnu_51_in_5, msg_to_check_it_11_cnu_52_in_0, msg_to_check_it_11_cnu_52_in_1, msg_to_check_it_11_cnu_52_in_2, msg_to_check_it_11_cnu_52_in_3, msg_to_check_it_11_cnu_52_in_4, msg_to_check_it_11_cnu_52_in_5, msg_to_check_it_11_cnu_53_in_0, msg_to_check_it_11_cnu_53_in_1, msg_to_check_it_11_cnu_53_in_2, msg_to_check_it_11_cnu_53_in_3, msg_to_check_it_11_cnu_53_in_4, msg_to_check_it_11_cnu_53_in_5, msg_to_check_it_11_cnu_54_in_0, msg_to_check_it_11_cnu_54_in_1, msg_to_check_it_11_cnu_54_in_2, msg_to_check_it_11_cnu_54_in_3, msg_to_check_it_11_cnu_54_in_4, msg_to_check_it_11_cnu_54_in_5, msg_to_check_it_11_cnu_55_in_0, msg_to_check_it_11_cnu_55_in_1, msg_to_check_it_11_cnu_55_in_2, msg_to_check_it_11_cnu_55_in_3, msg_to_check_it_11_cnu_55_in_4, msg_to_check_it_11_cnu_55_in_5, msg_to_check_it_11_cnu_56_in_0, msg_to_check_it_11_cnu_56_in_1, msg_to_check_it_11_cnu_56_in_2, msg_to_check_it_11_cnu_56_in_3, msg_to_check_it_11_cnu_56_in_4, msg_to_check_it_11_cnu_56_in_5, msg_to_check_it_11_cnu_57_in_0, msg_to_check_it_11_cnu_57_in_1, msg_to_check_it_11_cnu_57_in_2, msg_to_check_it_11_cnu_57_in_3, msg_to_check_it_11_cnu_57_in_4, msg_to_check_it_11_cnu_57_in_5, msg_to_check_it_11_cnu_58_in_0, msg_to_check_it_11_cnu_58_in_1, msg_to_check_it_11_cnu_58_in_2, msg_to_check_it_11_cnu_58_in_3, msg_to_check_it_11_cnu_58_in_4, msg_to_check_it_11_cnu_58_in_5, msg_to_check_it_11_cnu_59_in_0, msg_to_check_it_11_cnu_59_in_1, msg_to_check_it_11_cnu_59_in_2, msg_to_check_it_11_cnu_59_in_3, msg_to_check_it_11_cnu_59_in_4, msg_to_check_it_11_cnu_59_in_5, msg_to_check_it_11_cnu_60_in_0, msg_to_check_it_11_cnu_60_in_1, msg_to_check_it_11_cnu_60_in_2, msg_to_check_it_11_cnu_60_in_3, msg_to_check_it_11_cnu_60_in_4, msg_to_check_it_11_cnu_60_in_5, msg_to_check_it_11_cnu_61_in_0, msg_to_check_it_11_cnu_61_in_1, msg_to_check_it_11_cnu_61_in_2, msg_to_check_it_11_cnu_61_in_3, msg_to_check_it_11_cnu_61_in_4, msg_to_check_it_11_cnu_61_in_5, msg_to_check_it_11_cnu_62_in_0, msg_to_check_it_11_cnu_62_in_1, msg_to_check_it_11_cnu_62_in_2, msg_to_check_it_11_cnu_62_in_3, msg_to_check_it_11_cnu_62_in_4, msg_to_check_it_11_cnu_62_in_5, msg_to_check_it_11_cnu_63_in_0, msg_to_check_it_11_cnu_63_in_1, msg_to_check_it_11_cnu_63_in_2, msg_to_check_it_11_cnu_63_in_3, msg_to_check_it_11_cnu_63_in_4, msg_to_check_it_11_cnu_63_in_5, msg_to_check_it_11_cnu_64_in_0, msg_to_check_it_11_cnu_64_in_1, msg_to_check_it_11_cnu_64_in_2, msg_to_check_it_11_cnu_64_in_3, msg_to_check_it_11_cnu_64_in_4, msg_to_check_it_11_cnu_64_in_5, msg_to_check_it_11_cnu_65_in_0, msg_to_check_it_11_cnu_65_in_1, msg_to_check_it_11_cnu_65_in_2, msg_to_check_it_11_cnu_65_in_3, msg_to_check_it_11_cnu_65_in_4, msg_to_check_it_11_cnu_65_in_5, msg_to_check_it_11_cnu_66_in_0, msg_to_check_it_11_cnu_66_in_1, msg_to_check_it_11_cnu_66_in_2, msg_to_check_it_11_cnu_66_in_3, msg_to_check_it_11_cnu_66_in_4, msg_to_check_it_11_cnu_66_in_5, msg_to_check_it_11_cnu_67_in_0, msg_to_check_it_11_cnu_67_in_1, msg_to_check_it_11_cnu_67_in_2, msg_to_check_it_11_cnu_67_in_3, msg_to_check_it_11_cnu_67_in_4, msg_to_check_it_11_cnu_67_in_5, msg_to_check_it_11_cnu_68_in_0, msg_to_check_it_11_cnu_68_in_1, msg_to_check_it_11_cnu_68_in_2, msg_to_check_it_11_cnu_68_in_3, msg_to_check_it_11_cnu_68_in_4, msg_to_check_it_11_cnu_68_in_5, msg_to_check_it_11_cnu_69_in_0, msg_to_check_it_11_cnu_69_in_1, msg_to_check_it_11_cnu_69_in_2, msg_to_check_it_11_cnu_69_in_3, msg_to_check_it_11_cnu_69_in_4, msg_to_check_it_11_cnu_69_in_5, msg_to_check_it_11_cnu_70_in_0, msg_to_check_it_11_cnu_70_in_1, msg_to_check_it_11_cnu_70_in_2, msg_to_check_it_11_cnu_70_in_3, msg_to_check_it_11_cnu_70_in_4, msg_to_check_it_11_cnu_70_in_5, msg_to_check_it_11_cnu_71_in_0, msg_to_check_it_11_cnu_71_in_1, msg_to_check_it_11_cnu_71_in_2, msg_to_check_it_11_cnu_71_in_3, msg_to_check_it_11_cnu_71_in_4, msg_to_check_it_11_cnu_71_in_5, msg_to_check_it_11_cnu_72_in_0, msg_to_check_it_11_cnu_72_in_1, msg_to_check_it_11_cnu_72_in_2, msg_to_check_it_11_cnu_72_in_3, msg_to_check_it_11_cnu_72_in_4, msg_to_check_it_11_cnu_72_in_5, msg_to_check_it_11_cnu_73_in_0, msg_to_check_it_11_cnu_73_in_1, msg_to_check_it_11_cnu_73_in_2, msg_to_check_it_11_cnu_73_in_3, msg_to_check_it_11_cnu_73_in_4, msg_to_check_it_11_cnu_73_in_5, msg_to_check_it_11_cnu_74_in_0, msg_to_check_it_11_cnu_74_in_1, msg_to_check_it_11_cnu_74_in_2, msg_to_check_it_11_cnu_74_in_3, msg_to_check_it_11_cnu_74_in_4, msg_to_check_it_11_cnu_74_in_5, msg_to_check_it_11_cnu_75_in_0, msg_to_check_it_11_cnu_75_in_1, msg_to_check_it_11_cnu_75_in_2, msg_to_check_it_11_cnu_75_in_3, msg_to_check_it_11_cnu_75_in_4, msg_to_check_it_11_cnu_75_in_5, msg_to_check_it_11_cnu_76_in_0, msg_to_check_it_11_cnu_76_in_1, msg_to_check_it_11_cnu_76_in_2, msg_to_check_it_11_cnu_76_in_3, msg_to_check_it_11_cnu_76_in_4, msg_to_check_it_11_cnu_76_in_5, msg_to_check_it_11_cnu_77_in_0, msg_to_check_it_11_cnu_77_in_1, msg_to_check_it_11_cnu_77_in_2, msg_to_check_it_11_cnu_77_in_3, msg_to_check_it_11_cnu_77_in_4, msg_to_check_it_11_cnu_77_in_5, msg_to_check_it_11_cnu_78_in_0, msg_to_check_it_11_cnu_78_in_1, msg_to_check_it_11_cnu_78_in_2, msg_to_check_it_11_cnu_78_in_3, msg_to_check_it_11_cnu_78_in_4, msg_to_check_it_11_cnu_78_in_5, msg_to_check_it_11_cnu_79_in_0, msg_to_check_it_11_cnu_79_in_1, msg_to_check_it_11_cnu_79_in_2, msg_to_check_it_11_cnu_79_in_3, msg_to_check_it_11_cnu_79_in_4, msg_to_check_it_11_cnu_79_in_5, msg_to_check_it_11_cnu_80_in_0, msg_to_check_it_11_cnu_80_in_1, msg_to_check_it_11_cnu_80_in_2, msg_to_check_it_11_cnu_80_in_3, msg_to_check_it_11_cnu_80_in_4, msg_to_check_it_11_cnu_80_in_5, msg_to_check_it_11_cnu_81_in_0, msg_to_check_it_11_cnu_81_in_1, msg_to_check_it_11_cnu_81_in_2, msg_to_check_it_11_cnu_81_in_3, msg_to_check_it_11_cnu_81_in_4, msg_to_check_it_11_cnu_81_in_5, msg_to_check_it_11_cnu_82_in_0, msg_to_check_it_11_cnu_82_in_1, msg_to_check_it_11_cnu_82_in_2, msg_to_check_it_11_cnu_82_in_3, msg_to_check_it_11_cnu_82_in_4, msg_to_check_it_11_cnu_82_in_5, msg_to_check_it_11_cnu_83_in_0, msg_to_check_it_11_cnu_83_in_1, msg_to_check_it_11_cnu_83_in_2, msg_to_check_it_11_cnu_83_in_3, msg_to_check_it_11_cnu_83_in_4, msg_to_check_it_11_cnu_83_in_5, msg_to_check_it_11_cnu_84_in_0, msg_to_check_it_11_cnu_84_in_1, msg_to_check_it_11_cnu_84_in_2, msg_to_check_it_11_cnu_84_in_3, msg_to_check_it_11_cnu_84_in_4, msg_to_check_it_11_cnu_84_in_5, msg_to_check_it_11_cnu_85_in_0, msg_to_check_it_11_cnu_85_in_1, msg_to_check_it_11_cnu_85_in_2, msg_to_check_it_11_cnu_85_in_3, msg_to_check_it_11_cnu_85_in_4, msg_to_check_it_11_cnu_85_in_5, msg_to_check_it_11_cnu_86_in_0, msg_to_check_it_11_cnu_86_in_1, msg_to_check_it_11_cnu_86_in_2, msg_to_check_it_11_cnu_86_in_3, msg_to_check_it_11_cnu_86_in_4, msg_to_check_it_11_cnu_86_in_5, msg_to_check_it_11_cnu_87_in_0, msg_to_check_it_11_cnu_87_in_1, msg_to_check_it_11_cnu_87_in_2, msg_to_check_it_11_cnu_87_in_3, msg_to_check_it_11_cnu_87_in_4, msg_to_check_it_11_cnu_87_in_5, msg_to_check_it_11_cnu_88_in_0, msg_to_check_it_11_cnu_88_in_1, msg_to_check_it_11_cnu_88_in_2, msg_to_check_it_11_cnu_88_in_3, msg_to_check_it_11_cnu_88_in_4, msg_to_check_it_11_cnu_88_in_5, msg_to_check_it_11_cnu_89_in_0, msg_to_check_it_11_cnu_89_in_1, msg_to_check_it_11_cnu_89_in_2, msg_to_check_it_11_cnu_89_in_3, msg_to_check_it_11_cnu_89_in_4, msg_to_check_it_11_cnu_89_in_5, msg_to_check_it_11_cnu_90_in_0, msg_to_check_it_11_cnu_90_in_1, msg_to_check_it_11_cnu_90_in_2, msg_to_check_it_11_cnu_90_in_3, msg_to_check_it_11_cnu_90_in_4, msg_to_check_it_11_cnu_90_in_5, msg_to_check_it_11_cnu_91_in_0, msg_to_check_it_11_cnu_91_in_1, msg_to_check_it_11_cnu_91_in_2, msg_to_check_it_11_cnu_91_in_3, msg_to_check_it_11_cnu_91_in_4, msg_to_check_it_11_cnu_91_in_5, msg_to_check_it_11_cnu_92_in_0, msg_to_check_it_11_cnu_92_in_1, msg_to_check_it_11_cnu_92_in_2, msg_to_check_it_11_cnu_92_in_3, msg_to_check_it_11_cnu_92_in_4, msg_to_check_it_11_cnu_92_in_5, msg_to_check_it_11_cnu_93_in_0, msg_to_check_it_11_cnu_93_in_1, msg_to_check_it_11_cnu_93_in_2, msg_to_check_it_11_cnu_93_in_3, msg_to_check_it_11_cnu_93_in_4, msg_to_check_it_11_cnu_93_in_5, msg_to_check_it_11_cnu_94_in_0, msg_to_check_it_11_cnu_94_in_1, msg_to_check_it_11_cnu_94_in_2, msg_to_check_it_11_cnu_94_in_3, msg_to_check_it_11_cnu_94_in_4, msg_to_check_it_11_cnu_94_in_5, msg_to_check_it_11_cnu_95_in_0, msg_to_check_it_11_cnu_95_in_1, msg_to_check_it_11_cnu_95_in_2, msg_to_check_it_11_cnu_95_in_3, msg_to_check_it_11_cnu_95_in_4, msg_to_check_it_11_cnu_95_in_5, msg_to_check_it_11_cnu_96_in_0, msg_to_check_it_11_cnu_96_in_1, msg_to_check_it_11_cnu_96_in_2, msg_to_check_it_11_cnu_96_in_3, msg_to_check_it_11_cnu_96_in_4, msg_to_check_it_11_cnu_96_in_5, msg_to_check_it_11_cnu_97_in_0, msg_to_check_it_11_cnu_97_in_1, msg_to_check_it_11_cnu_97_in_2, msg_to_check_it_11_cnu_97_in_3, msg_to_check_it_11_cnu_97_in_4, msg_to_check_it_11_cnu_97_in_5, msg_to_check_it_11_cnu_98_in_0, msg_to_check_it_11_cnu_98_in_1, msg_to_check_it_11_cnu_98_in_2, msg_to_check_it_11_cnu_98_in_3, msg_to_check_it_11_cnu_98_in_4, msg_to_check_it_11_cnu_98_in_5, msg_to_check_it_12_cnu_0_in_0, msg_to_check_it_12_cnu_0_in_1, msg_to_check_it_12_cnu_0_in_2, msg_to_check_it_12_cnu_0_in_3, msg_to_check_it_12_cnu_0_in_4, msg_to_check_it_12_cnu_0_in_5, msg_to_check_it_12_cnu_1_in_0, msg_to_check_it_12_cnu_1_in_1, msg_to_check_it_12_cnu_1_in_2, msg_to_check_it_12_cnu_1_in_3, msg_to_check_it_12_cnu_1_in_4, msg_to_check_it_12_cnu_1_in_5, msg_to_check_it_12_cnu_2_in_0, msg_to_check_it_12_cnu_2_in_1, msg_to_check_it_12_cnu_2_in_2, msg_to_check_it_12_cnu_2_in_3, msg_to_check_it_12_cnu_2_in_4, msg_to_check_it_12_cnu_2_in_5, msg_to_check_it_12_cnu_3_in_0, msg_to_check_it_12_cnu_3_in_1, msg_to_check_it_12_cnu_3_in_2, msg_to_check_it_12_cnu_3_in_3, msg_to_check_it_12_cnu_3_in_4, msg_to_check_it_12_cnu_3_in_5, msg_to_check_it_12_cnu_4_in_0, msg_to_check_it_12_cnu_4_in_1, msg_to_check_it_12_cnu_4_in_2, msg_to_check_it_12_cnu_4_in_3, msg_to_check_it_12_cnu_4_in_4, msg_to_check_it_12_cnu_4_in_5, msg_to_check_it_12_cnu_5_in_0, msg_to_check_it_12_cnu_5_in_1, msg_to_check_it_12_cnu_5_in_2, msg_to_check_it_12_cnu_5_in_3, msg_to_check_it_12_cnu_5_in_4, msg_to_check_it_12_cnu_5_in_5, msg_to_check_it_12_cnu_6_in_0, msg_to_check_it_12_cnu_6_in_1, msg_to_check_it_12_cnu_6_in_2, msg_to_check_it_12_cnu_6_in_3, msg_to_check_it_12_cnu_6_in_4, msg_to_check_it_12_cnu_6_in_5, msg_to_check_it_12_cnu_7_in_0, msg_to_check_it_12_cnu_7_in_1, msg_to_check_it_12_cnu_7_in_2, msg_to_check_it_12_cnu_7_in_3, msg_to_check_it_12_cnu_7_in_4, msg_to_check_it_12_cnu_7_in_5, msg_to_check_it_12_cnu_8_in_0, msg_to_check_it_12_cnu_8_in_1, msg_to_check_it_12_cnu_8_in_2, msg_to_check_it_12_cnu_8_in_3, msg_to_check_it_12_cnu_8_in_4, msg_to_check_it_12_cnu_8_in_5, msg_to_check_it_12_cnu_9_in_0, msg_to_check_it_12_cnu_9_in_1, msg_to_check_it_12_cnu_9_in_2, msg_to_check_it_12_cnu_9_in_3, msg_to_check_it_12_cnu_9_in_4, msg_to_check_it_12_cnu_9_in_5, msg_to_check_it_12_cnu_10_in_0, msg_to_check_it_12_cnu_10_in_1, msg_to_check_it_12_cnu_10_in_2, msg_to_check_it_12_cnu_10_in_3, msg_to_check_it_12_cnu_10_in_4, msg_to_check_it_12_cnu_10_in_5, msg_to_check_it_12_cnu_11_in_0, msg_to_check_it_12_cnu_11_in_1, msg_to_check_it_12_cnu_11_in_2, msg_to_check_it_12_cnu_11_in_3, msg_to_check_it_12_cnu_11_in_4, msg_to_check_it_12_cnu_11_in_5, msg_to_check_it_12_cnu_12_in_0, msg_to_check_it_12_cnu_12_in_1, msg_to_check_it_12_cnu_12_in_2, msg_to_check_it_12_cnu_12_in_3, msg_to_check_it_12_cnu_12_in_4, msg_to_check_it_12_cnu_12_in_5, msg_to_check_it_12_cnu_13_in_0, msg_to_check_it_12_cnu_13_in_1, msg_to_check_it_12_cnu_13_in_2, msg_to_check_it_12_cnu_13_in_3, msg_to_check_it_12_cnu_13_in_4, msg_to_check_it_12_cnu_13_in_5, msg_to_check_it_12_cnu_14_in_0, msg_to_check_it_12_cnu_14_in_1, msg_to_check_it_12_cnu_14_in_2, msg_to_check_it_12_cnu_14_in_3, msg_to_check_it_12_cnu_14_in_4, msg_to_check_it_12_cnu_14_in_5, msg_to_check_it_12_cnu_15_in_0, msg_to_check_it_12_cnu_15_in_1, msg_to_check_it_12_cnu_15_in_2, msg_to_check_it_12_cnu_15_in_3, msg_to_check_it_12_cnu_15_in_4, msg_to_check_it_12_cnu_15_in_5, msg_to_check_it_12_cnu_16_in_0, msg_to_check_it_12_cnu_16_in_1, msg_to_check_it_12_cnu_16_in_2, msg_to_check_it_12_cnu_16_in_3, msg_to_check_it_12_cnu_16_in_4, msg_to_check_it_12_cnu_16_in_5, msg_to_check_it_12_cnu_17_in_0, msg_to_check_it_12_cnu_17_in_1, msg_to_check_it_12_cnu_17_in_2, msg_to_check_it_12_cnu_17_in_3, msg_to_check_it_12_cnu_17_in_4, msg_to_check_it_12_cnu_17_in_5, msg_to_check_it_12_cnu_18_in_0, msg_to_check_it_12_cnu_18_in_1, msg_to_check_it_12_cnu_18_in_2, msg_to_check_it_12_cnu_18_in_3, msg_to_check_it_12_cnu_18_in_4, msg_to_check_it_12_cnu_18_in_5, msg_to_check_it_12_cnu_19_in_0, msg_to_check_it_12_cnu_19_in_1, msg_to_check_it_12_cnu_19_in_2, msg_to_check_it_12_cnu_19_in_3, msg_to_check_it_12_cnu_19_in_4, msg_to_check_it_12_cnu_19_in_5, msg_to_check_it_12_cnu_20_in_0, msg_to_check_it_12_cnu_20_in_1, msg_to_check_it_12_cnu_20_in_2, msg_to_check_it_12_cnu_20_in_3, msg_to_check_it_12_cnu_20_in_4, msg_to_check_it_12_cnu_20_in_5, msg_to_check_it_12_cnu_21_in_0, msg_to_check_it_12_cnu_21_in_1, msg_to_check_it_12_cnu_21_in_2, msg_to_check_it_12_cnu_21_in_3, msg_to_check_it_12_cnu_21_in_4, msg_to_check_it_12_cnu_21_in_5, msg_to_check_it_12_cnu_22_in_0, msg_to_check_it_12_cnu_22_in_1, msg_to_check_it_12_cnu_22_in_2, msg_to_check_it_12_cnu_22_in_3, msg_to_check_it_12_cnu_22_in_4, msg_to_check_it_12_cnu_22_in_5, msg_to_check_it_12_cnu_23_in_0, msg_to_check_it_12_cnu_23_in_1, msg_to_check_it_12_cnu_23_in_2, msg_to_check_it_12_cnu_23_in_3, msg_to_check_it_12_cnu_23_in_4, msg_to_check_it_12_cnu_23_in_5, msg_to_check_it_12_cnu_24_in_0, msg_to_check_it_12_cnu_24_in_1, msg_to_check_it_12_cnu_24_in_2, msg_to_check_it_12_cnu_24_in_3, msg_to_check_it_12_cnu_24_in_4, msg_to_check_it_12_cnu_24_in_5, msg_to_check_it_12_cnu_25_in_0, msg_to_check_it_12_cnu_25_in_1, msg_to_check_it_12_cnu_25_in_2, msg_to_check_it_12_cnu_25_in_3, msg_to_check_it_12_cnu_25_in_4, msg_to_check_it_12_cnu_25_in_5, msg_to_check_it_12_cnu_26_in_0, msg_to_check_it_12_cnu_26_in_1, msg_to_check_it_12_cnu_26_in_2, msg_to_check_it_12_cnu_26_in_3, msg_to_check_it_12_cnu_26_in_4, msg_to_check_it_12_cnu_26_in_5, msg_to_check_it_12_cnu_27_in_0, msg_to_check_it_12_cnu_27_in_1, msg_to_check_it_12_cnu_27_in_2, msg_to_check_it_12_cnu_27_in_3, msg_to_check_it_12_cnu_27_in_4, msg_to_check_it_12_cnu_27_in_5, msg_to_check_it_12_cnu_28_in_0, msg_to_check_it_12_cnu_28_in_1, msg_to_check_it_12_cnu_28_in_2, msg_to_check_it_12_cnu_28_in_3, msg_to_check_it_12_cnu_28_in_4, msg_to_check_it_12_cnu_28_in_5, msg_to_check_it_12_cnu_29_in_0, msg_to_check_it_12_cnu_29_in_1, msg_to_check_it_12_cnu_29_in_2, msg_to_check_it_12_cnu_29_in_3, msg_to_check_it_12_cnu_29_in_4, msg_to_check_it_12_cnu_29_in_5, msg_to_check_it_12_cnu_30_in_0, msg_to_check_it_12_cnu_30_in_1, msg_to_check_it_12_cnu_30_in_2, msg_to_check_it_12_cnu_30_in_3, msg_to_check_it_12_cnu_30_in_4, msg_to_check_it_12_cnu_30_in_5, msg_to_check_it_12_cnu_31_in_0, msg_to_check_it_12_cnu_31_in_1, msg_to_check_it_12_cnu_31_in_2, msg_to_check_it_12_cnu_31_in_3, msg_to_check_it_12_cnu_31_in_4, msg_to_check_it_12_cnu_31_in_5, msg_to_check_it_12_cnu_32_in_0, msg_to_check_it_12_cnu_32_in_1, msg_to_check_it_12_cnu_32_in_2, msg_to_check_it_12_cnu_32_in_3, msg_to_check_it_12_cnu_32_in_4, msg_to_check_it_12_cnu_32_in_5, msg_to_check_it_12_cnu_33_in_0, msg_to_check_it_12_cnu_33_in_1, msg_to_check_it_12_cnu_33_in_2, msg_to_check_it_12_cnu_33_in_3, msg_to_check_it_12_cnu_33_in_4, msg_to_check_it_12_cnu_33_in_5, msg_to_check_it_12_cnu_34_in_0, msg_to_check_it_12_cnu_34_in_1, msg_to_check_it_12_cnu_34_in_2, msg_to_check_it_12_cnu_34_in_3, msg_to_check_it_12_cnu_34_in_4, msg_to_check_it_12_cnu_34_in_5, msg_to_check_it_12_cnu_35_in_0, msg_to_check_it_12_cnu_35_in_1, msg_to_check_it_12_cnu_35_in_2, msg_to_check_it_12_cnu_35_in_3, msg_to_check_it_12_cnu_35_in_4, msg_to_check_it_12_cnu_35_in_5, msg_to_check_it_12_cnu_36_in_0, msg_to_check_it_12_cnu_36_in_1, msg_to_check_it_12_cnu_36_in_2, msg_to_check_it_12_cnu_36_in_3, msg_to_check_it_12_cnu_36_in_4, msg_to_check_it_12_cnu_36_in_5, msg_to_check_it_12_cnu_37_in_0, msg_to_check_it_12_cnu_37_in_1, msg_to_check_it_12_cnu_37_in_2, msg_to_check_it_12_cnu_37_in_3, msg_to_check_it_12_cnu_37_in_4, msg_to_check_it_12_cnu_37_in_5, msg_to_check_it_12_cnu_38_in_0, msg_to_check_it_12_cnu_38_in_1, msg_to_check_it_12_cnu_38_in_2, msg_to_check_it_12_cnu_38_in_3, msg_to_check_it_12_cnu_38_in_4, msg_to_check_it_12_cnu_38_in_5, msg_to_check_it_12_cnu_39_in_0, msg_to_check_it_12_cnu_39_in_1, msg_to_check_it_12_cnu_39_in_2, msg_to_check_it_12_cnu_39_in_3, msg_to_check_it_12_cnu_39_in_4, msg_to_check_it_12_cnu_39_in_5, msg_to_check_it_12_cnu_40_in_0, msg_to_check_it_12_cnu_40_in_1, msg_to_check_it_12_cnu_40_in_2, msg_to_check_it_12_cnu_40_in_3, msg_to_check_it_12_cnu_40_in_4, msg_to_check_it_12_cnu_40_in_5, msg_to_check_it_12_cnu_41_in_0, msg_to_check_it_12_cnu_41_in_1, msg_to_check_it_12_cnu_41_in_2, msg_to_check_it_12_cnu_41_in_3, msg_to_check_it_12_cnu_41_in_4, msg_to_check_it_12_cnu_41_in_5, msg_to_check_it_12_cnu_42_in_0, msg_to_check_it_12_cnu_42_in_1, msg_to_check_it_12_cnu_42_in_2, msg_to_check_it_12_cnu_42_in_3, msg_to_check_it_12_cnu_42_in_4, msg_to_check_it_12_cnu_42_in_5, msg_to_check_it_12_cnu_43_in_0, msg_to_check_it_12_cnu_43_in_1, msg_to_check_it_12_cnu_43_in_2, msg_to_check_it_12_cnu_43_in_3, msg_to_check_it_12_cnu_43_in_4, msg_to_check_it_12_cnu_43_in_5, msg_to_check_it_12_cnu_44_in_0, msg_to_check_it_12_cnu_44_in_1, msg_to_check_it_12_cnu_44_in_2, msg_to_check_it_12_cnu_44_in_3, msg_to_check_it_12_cnu_44_in_4, msg_to_check_it_12_cnu_44_in_5, msg_to_check_it_12_cnu_45_in_0, msg_to_check_it_12_cnu_45_in_1, msg_to_check_it_12_cnu_45_in_2, msg_to_check_it_12_cnu_45_in_3, msg_to_check_it_12_cnu_45_in_4, msg_to_check_it_12_cnu_45_in_5, msg_to_check_it_12_cnu_46_in_0, msg_to_check_it_12_cnu_46_in_1, msg_to_check_it_12_cnu_46_in_2, msg_to_check_it_12_cnu_46_in_3, msg_to_check_it_12_cnu_46_in_4, msg_to_check_it_12_cnu_46_in_5, msg_to_check_it_12_cnu_47_in_0, msg_to_check_it_12_cnu_47_in_1, msg_to_check_it_12_cnu_47_in_2, msg_to_check_it_12_cnu_47_in_3, msg_to_check_it_12_cnu_47_in_4, msg_to_check_it_12_cnu_47_in_5, msg_to_check_it_12_cnu_48_in_0, msg_to_check_it_12_cnu_48_in_1, msg_to_check_it_12_cnu_48_in_2, msg_to_check_it_12_cnu_48_in_3, msg_to_check_it_12_cnu_48_in_4, msg_to_check_it_12_cnu_48_in_5, msg_to_check_it_12_cnu_49_in_0, msg_to_check_it_12_cnu_49_in_1, msg_to_check_it_12_cnu_49_in_2, msg_to_check_it_12_cnu_49_in_3, msg_to_check_it_12_cnu_49_in_4, msg_to_check_it_12_cnu_49_in_5, msg_to_check_it_12_cnu_50_in_0, msg_to_check_it_12_cnu_50_in_1, msg_to_check_it_12_cnu_50_in_2, msg_to_check_it_12_cnu_50_in_3, msg_to_check_it_12_cnu_50_in_4, msg_to_check_it_12_cnu_50_in_5, msg_to_check_it_12_cnu_51_in_0, msg_to_check_it_12_cnu_51_in_1, msg_to_check_it_12_cnu_51_in_2, msg_to_check_it_12_cnu_51_in_3, msg_to_check_it_12_cnu_51_in_4, msg_to_check_it_12_cnu_51_in_5, msg_to_check_it_12_cnu_52_in_0, msg_to_check_it_12_cnu_52_in_1, msg_to_check_it_12_cnu_52_in_2, msg_to_check_it_12_cnu_52_in_3, msg_to_check_it_12_cnu_52_in_4, msg_to_check_it_12_cnu_52_in_5, msg_to_check_it_12_cnu_53_in_0, msg_to_check_it_12_cnu_53_in_1, msg_to_check_it_12_cnu_53_in_2, msg_to_check_it_12_cnu_53_in_3, msg_to_check_it_12_cnu_53_in_4, msg_to_check_it_12_cnu_53_in_5, msg_to_check_it_12_cnu_54_in_0, msg_to_check_it_12_cnu_54_in_1, msg_to_check_it_12_cnu_54_in_2, msg_to_check_it_12_cnu_54_in_3, msg_to_check_it_12_cnu_54_in_4, msg_to_check_it_12_cnu_54_in_5, msg_to_check_it_12_cnu_55_in_0, msg_to_check_it_12_cnu_55_in_1, msg_to_check_it_12_cnu_55_in_2, msg_to_check_it_12_cnu_55_in_3, msg_to_check_it_12_cnu_55_in_4, msg_to_check_it_12_cnu_55_in_5, msg_to_check_it_12_cnu_56_in_0, msg_to_check_it_12_cnu_56_in_1, msg_to_check_it_12_cnu_56_in_2, msg_to_check_it_12_cnu_56_in_3, msg_to_check_it_12_cnu_56_in_4, msg_to_check_it_12_cnu_56_in_5, msg_to_check_it_12_cnu_57_in_0, msg_to_check_it_12_cnu_57_in_1, msg_to_check_it_12_cnu_57_in_2, msg_to_check_it_12_cnu_57_in_3, msg_to_check_it_12_cnu_57_in_4, msg_to_check_it_12_cnu_57_in_5, msg_to_check_it_12_cnu_58_in_0, msg_to_check_it_12_cnu_58_in_1, msg_to_check_it_12_cnu_58_in_2, msg_to_check_it_12_cnu_58_in_3, msg_to_check_it_12_cnu_58_in_4, msg_to_check_it_12_cnu_58_in_5, msg_to_check_it_12_cnu_59_in_0, msg_to_check_it_12_cnu_59_in_1, msg_to_check_it_12_cnu_59_in_2, msg_to_check_it_12_cnu_59_in_3, msg_to_check_it_12_cnu_59_in_4, msg_to_check_it_12_cnu_59_in_5, msg_to_check_it_12_cnu_60_in_0, msg_to_check_it_12_cnu_60_in_1, msg_to_check_it_12_cnu_60_in_2, msg_to_check_it_12_cnu_60_in_3, msg_to_check_it_12_cnu_60_in_4, msg_to_check_it_12_cnu_60_in_5, msg_to_check_it_12_cnu_61_in_0, msg_to_check_it_12_cnu_61_in_1, msg_to_check_it_12_cnu_61_in_2, msg_to_check_it_12_cnu_61_in_3, msg_to_check_it_12_cnu_61_in_4, msg_to_check_it_12_cnu_61_in_5, msg_to_check_it_12_cnu_62_in_0, msg_to_check_it_12_cnu_62_in_1, msg_to_check_it_12_cnu_62_in_2, msg_to_check_it_12_cnu_62_in_3, msg_to_check_it_12_cnu_62_in_4, msg_to_check_it_12_cnu_62_in_5, msg_to_check_it_12_cnu_63_in_0, msg_to_check_it_12_cnu_63_in_1, msg_to_check_it_12_cnu_63_in_2, msg_to_check_it_12_cnu_63_in_3, msg_to_check_it_12_cnu_63_in_4, msg_to_check_it_12_cnu_63_in_5, msg_to_check_it_12_cnu_64_in_0, msg_to_check_it_12_cnu_64_in_1, msg_to_check_it_12_cnu_64_in_2, msg_to_check_it_12_cnu_64_in_3, msg_to_check_it_12_cnu_64_in_4, msg_to_check_it_12_cnu_64_in_5, msg_to_check_it_12_cnu_65_in_0, msg_to_check_it_12_cnu_65_in_1, msg_to_check_it_12_cnu_65_in_2, msg_to_check_it_12_cnu_65_in_3, msg_to_check_it_12_cnu_65_in_4, msg_to_check_it_12_cnu_65_in_5, msg_to_check_it_12_cnu_66_in_0, msg_to_check_it_12_cnu_66_in_1, msg_to_check_it_12_cnu_66_in_2, msg_to_check_it_12_cnu_66_in_3, msg_to_check_it_12_cnu_66_in_4, msg_to_check_it_12_cnu_66_in_5, msg_to_check_it_12_cnu_67_in_0, msg_to_check_it_12_cnu_67_in_1, msg_to_check_it_12_cnu_67_in_2, msg_to_check_it_12_cnu_67_in_3, msg_to_check_it_12_cnu_67_in_4, msg_to_check_it_12_cnu_67_in_5, msg_to_check_it_12_cnu_68_in_0, msg_to_check_it_12_cnu_68_in_1, msg_to_check_it_12_cnu_68_in_2, msg_to_check_it_12_cnu_68_in_3, msg_to_check_it_12_cnu_68_in_4, msg_to_check_it_12_cnu_68_in_5, msg_to_check_it_12_cnu_69_in_0, msg_to_check_it_12_cnu_69_in_1, msg_to_check_it_12_cnu_69_in_2, msg_to_check_it_12_cnu_69_in_3, msg_to_check_it_12_cnu_69_in_4, msg_to_check_it_12_cnu_69_in_5, msg_to_check_it_12_cnu_70_in_0, msg_to_check_it_12_cnu_70_in_1, msg_to_check_it_12_cnu_70_in_2, msg_to_check_it_12_cnu_70_in_3, msg_to_check_it_12_cnu_70_in_4, msg_to_check_it_12_cnu_70_in_5, msg_to_check_it_12_cnu_71_in_0, msg_to_check_it_12_cnu_71_in_1, msg_to_check_it_12_cnu_71_in_2, msg_to_check_it_12_cnu_71_in_3, msg_to_check_it_12_cnu_71_in_4, msg_to_check_it_12_cnu_71_in_5, msg_to_check_it_12_cnu_72_in_0, msg_to_check_it_12_cnu_72_in_1, msg_to_check_it_12_cnu_72_in_2, msg_to_check_it_12_cnu_72_in_3, msg_to_check_it_12_cnu_72_in_4, msg_to_check_it_12_cnu_72_in_5, msg_to_check_it_12_cnu_73_in_0, msg_to_check_it_12_cnu_73_in_1, msg_to_check_it_12_cnu_73_in_2, msg_to_check_it_12_cnu_73_in_3, msg_to_check_it_12_cnu_73_in_4, msg_to_check_it_12_cnu_73_in_5, msg_to_check_it_12_cnu_74_in_0, msg_to_check_it_12_cnu_74_in_1, msg_to_check_it_12_cnu_74_in_2, msg_to_check_it_12_cnu_74_in_3, msg_to_check_it_12_cnu_74_in_4, msg_to_check_it_12_cnu_74_in_5, msg_to_check_it_12_cnu_75_in_0, msg_to_check_it_12_cnu_75_in_1, msg_to_check_it_12_cnu_75_in_2, msg_to_check_it_12_cnu_75_in_3, msg_to_check_it_12_cnu_75_in_4, msg_to_check_it_12_cnu_75_in_5, msg_to_check_it_12_cnu_76_in_0, msg_to_check_it_12_cnu_76_in_1, msg_to_check_it_12_cnu_76_in_2, msg_to_check_it_12_cnu_76_in_3, msg_to_check_it_12_cnu_76_in_4, msg_to_check_it_12_cnu_76_in_5, msg_to_check_it_12_cnu_77_in_0, msg_to_check_it_12_cnu_77_in_1, msg_to_check_it_12_cnu_77_in_2, msg_to_check_it_12_cnu_77_in_3, msg_to_check_it_12_cnu_77_in_4, msg_to_check_it_12_cnu_77_in_5, msg_to_check_it_12_cnu_78_in_0, msg_to_check_it_12_cnu_78_in_1, msg_to_check_it_12_cnu_78_in_2, msg_to_check_it_12_cnu_78_in_3, msg_to_check_it_12_cnu_78_in_4, msg_to_check_it_12_cnu_78_in_5, msg_to_check_it_12_cnu_79_in_0, msg_to_check_it_12_cnu_79_in_1, msg_to_check_it_12_cnu_79_in_2, msg_to_check_it_12_cnu_79_in_3, msg_to_check_it_12_cnu_79_in_4, msg_to_check_it_12_cnu_79_in_5, msg_to_check_it_12_cnu_80_in_0, msg_to_check_it_12_cnu_80_in_1, msg_to_check_it_12_cnu_80_in_2, msg_to_check_it_12_cnu_80_in_3, msg_to_check_it_12_cnu_80_in_4, msg_to_check_it_12_cnu_80_in_5, msg_to_check_it_12_cnu_81_in_0, msg_to_check_it_12_cnu_81_in_1, msg_to_check_it_12_cnu_81_in_2, msg_to_check_it_12_cnu_81_in_3, msg_to_check_it_12_cnu_81_in_4, msg_to_check_it_12_cnu_81_in_5, msg_to_check_it_12_cnu_82_in_0, msg_to_check_it_12_cnu_82_in_1, msg_to_check_it_12_cnu_82_in_2, msg_to_check_it_12_cnu_82_in_3, msg_to_check_it_12_cnu_82_in_4, msg_to_check_it_12_cnu_82_in_5, msg_to_check_it_12_cnu_83_in_0, msg_to_check_it_12_cnu_83_in_1, msg_to_check_it_12_cnu_83_in_2, msg_to_check_it_12_cnu_83_in_3, msg_to_check_it_12_cnu_83_in_4, msg_to_check_it_12_cnu_83_in_5, msg_to_check_it_12_cnu_84_in_0, msg_to_check_it_12_cnu_84_in_1, msg_to_check_it_12_cnu_84_in_2, msg_to_check_it_12_cnu_84_in_3, msg_to_check_it_12_cnu_84_in_4, msg_to_check_it_12_cnu_84_in_5, msg_to_check_it_12_cnu_85_in_0, msg_to_check_it_12_cnu_85_in_1, msg_to_check_it_12_cnu_85_in_2, msg_to_check_it_12_cnu_85_in_3, msg_to_check_it_12_cnu_85_in_4, msg_to_check_it_12_cnu_85_in_5, msg_to_check_it_12_cnu_86_in_0, msg_to_check_it_12_cnu_86_in_1, msg_to_check_it_12_cnu_86_in_2, msg_to_check_it_12_cnu_86_in_3, msg_to_check_it_12_cnu_86_in_4, msg_to_check_it_12_cnu_86_in_5, msg_to_check_it_12_cnu_87_in_0, msg_to_check_it_12_cnu_87_in_1, msg_to_check_it_12_cnu_87_in_2, msg_to_check_it_12_cnu_87_in_3, msg_to_check_it_12_cnu_87_in_4, msg_to_check_it_12_cnu_87_in_5, msg_to_check_it_12_cnu_88_in_0, msg_to_check_it_12_cnu_88_in_1, msg_to_check_it_12_cnu_88_in_2, msg_to_check_it_12_cnu_88_in_3, msg_to_check_it_12_cnu_88_in_4, msg_to_check_it_12_cnu_88_in_5, msg_to_check_it_12_cnu_89_in_0, msg_to_check_it_12_cnu_89_in_1, msg_to_check_it_12_cnu_89_in_2, msg_to_check_it_12_cnu_89_in_3, msg_to_check_it_12_cnu_89_in_4, msg_to_check_it_12_cnu_89_in_5, msg_to_check_it_12_cnu_90_in_0, msg_to_check_it_12_cnu_90_in_1, msg_to_check_it_12_cnu_90_in_2, msg_to_check_it_12_cnu_90_in_3, msg_to_check_it_12_cnu_90_in_4, msg_to_check_it_12_cnu_90_in_5, msg_to_check_it_12_cnu_91_in_0, msg_to_check_it_12_cnu_91_in_1, msg_to_check_it_12_cnu_91_in_2, msg_to_check_it_12_cnu_91_in_3, msg_to_check_it_12_cnu_91_in_4, msg_to_check_it_12_cnu_91_in_5, msg_to_check_it_12_cnu_92_in_0, msg_to_check_it_12_cnu_92_in_1, msg_to_check_it_12_cnu_92_in_2, msg_to_check_it_12_cnu_92_in_3, msg_to_check_it_12_cnu_92_in_4, msg_to_check_it_12_cnu_92_in_5, msg_to_check_it_12_cnu_93_in_0, msg_to_check_it_12_cnu_93_in_1, msg_to_check_it_12_cnu_93_in_2, msg_to_check_it_12_cnu_93_in_3, msg_to_check_it_12_cnu_93_in_4, msg_to_check_it_12_cnu_93_in_5, msg_to_check_it_12_cnu_94_in_0, msg_to_check_it_12_cnu_94_in_1, msg_to_check_it_12_cnu_94_in_2, msg_to_check_it_12_cnu_94_in_3, msg_to_check_it_12_cnu_94_in_4, msg_to_check_it_12_cnu_94_in_5, msg_to_check_it_12_cnu_95_in_0, msg_to_check_it_12_cnu_95_in_1, msg_to_check_it_12_cnu_95_in_2, msg_to_check_it_12_cnu_95_in_3, msg_to_check_it_12_cnu_95_in_4, msg_to_check_it_12_cnu_95_in_5, msg_to_check_it_12_cnu_96_in_0, msg_to_check_it_12_cnu_96_in_1, msg_to_check_it_12_cnu_96_in_2, msg_to_check_it_12_cnu_96_in_3, msg_to_check_it_12_cnu_96_in_4, msg_to_check_it_12_cnu_96_in_5, msg_to_check_it_12_cnu_97_in_0, msg_to_check_it_12_cnu_97_in_1, msg_to_check_it_12_cnu_97_in_2, msg_to_check_it_12_cnu_97_in_3, msg_to_check_it_12_cnu_97_in_4, msg_to_check_it_12_cnu_97_in_5, msg_to_check_it_12_cnu_98_in_0, msg_to_check_it_12_cnu_98_in_1, msg_to_check_it_12_cnu_98_in_2, msg_to_check_it_12_cnu_98_in_3, msg_to_check_it_12_cnu_98_in_4, msg_to_check_it_12_cnu_98_in_5, msg_to_check_it_13_cnu_0_in_0, msg_to_check_it_13_cnu_0_in_1, msg_to_check_it_13_cnu_0_in_2, msg_to_check_it_13_cnu_0_in_3, msg_to_check_it_13_cnu_0_in_4, msg_to_check_it_13_cnu_0_in_5, msg_to_check_it_13_cnu_1_in_0, msg_to_check_it_13_cnu_1_in_1, msg_to_check_it_13_cnu_1_in_2, msg_to_check_it_13_cnu_1_in_3, msg_to_check_it_13_cnu_1_in_4, msg_to_check_it_13_cnu_1_in_5, msg_to_check_it_13_cnu_2_in_0, msg_to_check_it_13_cnu_2_in_1, msg_to_check_it_13_cnu_2_in_2, msg_to_check_it_13_cnu_2_in_3, msg_to_check_it_13_cnu_2_in_4, msg_to_check_it_13_cnu_2_in_5, msg_to_check_it_13_cnu_3_in_0, msg_to_check_it_13_cnu_3_in_1, msg_to_check_it_13_cnu_3_in_2, msg_to_check_it_13_cnu_3_in_3, msg_to_check_it_13_cnu_3_in_4, msg_to_check_it_13_cnu_3_in_5, msg_to_check_it_13_cnu_4_in_0, msg_to_check_it_13_cnu_4_in_1, msg_to_check_it_13_cnu_4_in_2, msg_to_check_it_13_cnu_4_in_3, msg_to_check_it_13_cnu_4_in_4, msg_to_check_it_13_cnu_4_in_5, msg_to_check_it_13_cnu_5_in_0, msg_to_check_it_13_cnu_5_in_1, msg_to_check_it_13_cnu_5_in_2, msg_to_check_it_13_cnu_5_in_3, msg_to_check_it_13_cnu_5_in_4, msg_to_check_it_13_cnu_5_in_5, msg_to_check_it_13_cnu_6_in_0, msg_to_check_it_13_cnu_6_in_1, msg_to_check_it_13_cnu_6_in_2, msg_to_check_it_13_cnu_6_in_3, msg_to_check_it_13_cnu_6_in_4, msg_to_check_it_13_cnu_6_in_5, msg_to_check_it_13_cnu_7_in_0, msg_to_check_it_13_cnu_7_in_1, msg_to_check_it_13_cnu_7_in_2, msg_to_check_it_13_cnu_7_in_3, msg_to_check_it_13_cnu_7_in_4, msg_to_check_it_13_cnu_7_in_5, msg_to_check_it_13_cnu_8_in_0, msg_to_check_it_13_cnu_8_in_1, msg_to_check_it_13_cnu_8_in_2, msg_to_check_it_13_cnu_8_in_3, msg_to_check_it_13_cnu_8_in_4, msg_to_check_it_13_cnu_8_in_5, msg_to_check_it_13_cnu_9_in_0, msg_to_check_it_13_cnu_9_in_1, msg_to_check_it_13_cnu_9_in_2, msg_to_check_it_13_cnu_9_in_3, msg_to_check_it_13_cnu_9_in_4, msg_to_check_it_13_cnu_9_in_5, msg_to_check_it_13_cnu_10_in_0, msg_to_check_it_13_cnu_10_in_1, msg_to_check_it_13_cnu_10_in_2, msg_to_check_it_13_cnu_10_in_3, msg_to_check_it_13_cnu_10_in_4, msg_to_check_it_13_cnu_10_in_5, msg_to_check_it_13_cnu_11_in_0, msg_to_check_it_13_cnu_11_in_1, msg_to_check_it_13_cnu_11_in_2, msg_to_check_it_13_cnu_11_in_3, msg_to_check_it_13_cnu_11_in_4, msg_to_check_it_13_cnu_11_in_5, msg_to_check_it_13_cnu_12_in_0, msg_to_check_it_13_cnu_12_in_1, msg_to_check_it_13_cnu_12_in_2, msg_to_check_it_13_cnu_12_in_3, msg_to_check_it_13_cnu_12_in_4, msg_to_check_it_13_cnu_12_in_5, msg_to_check_it_13_cnu_13_in_0, msg_to_check_it_13_cnu_13_in_1, msg_to_check_it_13_cnu_13_in_2, msg_to_check_it_13_cnu_13_in_3, msg_to_check_it_13_cnu_13_in_4, msg_to_check_it_13_cnu_13_in_5, msg_to_check_it_13_cnu_14_in_0, msg_to_check_it_13_cnu_14_in_1, msg_to_check_it_13_cnu_14_in_2, msg_to_check_it_13_cnu_14_in_3, msg_to_check_it_13_cnu_14_in_4, msg_to_check_it_13_cnu_14_in_5, msg_to_check_it_13_cnu_15_in_0, msg_to_check_it_13_cnu_15_in_1, msg_to_check_it_13_cnu_15_in_2, msg_to_check_it_13_cnu_15_in_3, msg_to_check_it_13_cnu_15_in_4, msg_to_check_it_13_cnu_15_in_5, msg_to_check_it_13_cnu_16_in_0, msg_to_check_it_13_cnu_16_in_1, msg_to_check_it_13_cnu_16_in_2, msg_to_check_it_13_cnu_16_in_3, msg_to_check_it_13_cnu_16_in_4, msg_to_check_it_13_cnu_16_in_5, msg_to_check_it_13_cnu_17_in_0, msg_to_check_it_13_cnu_17_in_1, msg_to_check_it_13_cnu_17_in_2, msg_to_check_it_13_cnu_17_in_3, msg_to_check_it_13_cnu_17_in_4, msg_to_check_it_13_cnu_17_in_5, msg_to_check_it_13_cnu_18_in_0, msg_to_check_it_13_cnu_18_in_1, msg_to_check_it_13_cnu_18_in_2, msg_to_check_it_13_cnu_18_in_3, msg_to_check_it_13_cnu_18_in_4, msg_to_check_it_13_cnu_18_in_5, msg_to_check_it_13_cnu_19_in_0, msg_to_check_it_13_cnu_19_in_1, msg_to_check_it_13_cnu_19_in_2, msg_to_check_it_13_cnu_19_in_3, msg_to_check_it_13_cnu_19_in_4, msg_to_check_it_13_cnu_19_in_5, msg_to_check_it_13_cnu_20_in_0, msg_to_check_it_13_cnu_20_in_1, msg_to_check_it_13_cnu_20_in_2, msg_to_check_it_13_cnu_20_in_3, msg_to_check_it_13_cnu_20_in_4, msg_to_check_it_13_cnu_20_in_5, msg_to_check_it_13_cnu_21_in_0, msg_to_check_it_13_cnu_21_in_1, msg_to_check_it_13_cnu_21_in_2, msg_to_check_it_13_cnu_21_in_3, msg_to_check_it_13_cnu_21_in_4, msg_to_check_it_13_cnu_21_in_5, msg_to_check_it_13_cnu_22_in_0, msg_to_check_it_13_cnu_22_in_1, msg_to_check_it_13_cnu_22_in_2, msg_to_check_it_13_cnu_22_in_3, msg_to_check_it_13_cnu_22_in_4, msg_to_check_it_13_cnu_22_in_5, msg_to_check_it_13_cnu_23_in_0, msg_to_check_it_13_cnu_23_in_1, msg_to_check_it_13_cnu_23_in_2, msg_to_check_it_13_cnu_23_in_3, msg_to_check_it_13_cnu_23_in_4, msg_to_check_it_13_cnu_23_in_5, msg_to_check_it_13_cnu_24_in_0, msg_to_check_it_13_cnu_24_in_1, msg_to_check_it_13_cnu_24_in_2, msg_to_check_it_13_cnu_24_in_3, msg_to_check_it_13_cnu_24_in_4, msg_to_check_it_13_cnu_24_in_5, msg_to_check_it_13_cnu_25_in_0, msg_to_check_it_13_cnu_25_in_1, msg_to_check_it_13_cnu_25_in_2, msg_to_check_it_13_cnu_25_in_3, msg_to_check_it_13_cnu_25_in_4, msg_to_check_it_13_cnu_25_in_5, msg_to_check_it_13_cnu_26_in_0, msg_to_check_it_13_cnu_26_in_1, msg_to_check_it_13_cnu_26_in_2, msg_to_check_it_13_cnu_26_in_3, msg_to_check_it_13_cnu_26_in_4, msg_to_check_it_13_cnu_26_in_5, msg_to_check_it_13_cnu_27_in_0, msg_to_check_it_13_cnu_27_in_1, msg_to_check_it_13_cnu_27_in_2, msg_to_check_it_13_cnu_27_in_3, msg_to_check_it_13_cnu_27_in_4, msg_to_check_it_13_cnu_27_in_5, msg_to_check_it_13_cnu_28_in_0, msg_to_check_it_13_cnu_28_in_1, msg_to_check_it_13_cnu_28_in_2, msg_to_check_it_13_cnu_28_in_3, msg_to_check_it_13_cnu_28_in_4, msg_to_check_it_13_cnu_28_in_5, msg_to_check_it_13_cnu_29_in_0, msg_to_check_it_13_cnu_29_in_1, msg_to_check_it_13_cnu_29_in_2, msg_to_check_it_13_cnu_29_in_3, msg_to_check_it_13_cnu_29_in_4, msg_to_check_it_13_cnu_29_in_5, msg_to_check_it_13_cnu_30_in_0, msg_to_check_it_13_cnu_30_in_1, msg_to_check_it_13_cnu_30_in_2, msg_to_check_it_13_cnu_30_in_3, msg_to_check_it_13_cnu_30_in_4, msg_to_check_it_13_cnu_30_in_5, msg_to_check_it_13_cnu_31_in_0, msg_to_check_it_13_cnu_31_in_1, msg_to_check_it_13_cnu_31_in_2, msg_to_check_it_13_cnu_31_in_3, msg_to_check_it_13_cnu_31_in_4, msg_to_check_it_13_cnu_31_in_5, msg_to_check_it_13_cnu_32_in_0, msg_to_check_it_13_cnu_32_in_1, msg_to_check_it_13_cnu_32_in_2, msg_to_check_it_13_cnu_32_in_3, msg_to_check_it_13_cnu_32_in_4, msg_to_check_it_13_cnu_32_in_5, msg_to_check_it_13_cnu_33_in_0, msg_to_check_it_13_cnu_33_in_1, msg_to_check_it_13_cnu_33_in_2, msg_to_check_it_13_cnu_33_in_3, msg_to_check_it_13_cnu_33_in_4, msg_to_check_it_13_cnu_33_in_5, msg_to_check_it_13_cnu_34_in_0, msg_to_check_it_13_cnu_34_in_1, msg_to_check_it_13_cnu_34_in_2, msg_to_check_it_13_cnu_34_in_3, msg_to_check_it_13_cnu_34_in_4, msg_to_check_it_13_cnu_34_in_5, msg_to_check_it_13_cnu_35_in_0, msg_to_check_it_13_cnu_35_in_1, msg_to_check_it_13_cnu_35_in_2, msg_to_check_it_13_cnu_35_in_3, msg_to_check_it_13_cnu_35_in_4, msg_to_check_it_13_cnu_35_in_5, msg_to_check_it_13_cnu_36_in_0, msg_to_check_it_13_cnu_36_in_1, msg_to_check_it_13_cnu_36_in_2, msg_to_check_it_13_cnu_36_in_3, msg_to_check_it_13_cnu_36_in_4, msg_to_check_it_13_cnu_36_in_5, msg_to_check_it_13_cnu_37_in_0, msg_to_check_it_13_cnu_37_in_1, msg_to_check_it_13_cnu_37_in_2, msg_to_check_it_13_cnu_37_in_3, msg_to_check_it_13_cnu_37_in_4, msg_to_check_it_13_cnu_37_in_5, msg_to_check_it_13_cnu_38_in_0, msg_to_check_it_13_cnu_38_in_1, msg_to_check_it_13_cnu_38_in_2, msg_to_check_it_13_cnu_38_in_3, msg_to_check_it_13_cnu_38_in_4, msg_to_check_it_13_cnu_38_in_5, msg_to_check_it_13_cnu_39_in_0, msg_to_check_it_13_cnu_39_in_1, msg_to_check_it_13_cnu_39_in_2, msg_to_check_it_13_cnu_39_in_3, msg_to_check_it_13_cnu_39_in_4, msg_to_check_it_13_cnu_39_in_5, msg_to_check_it_13_cnu_40_in_0, msg_to_check_it_13_cnu_40_in_1, msg_to_check_it_13_cnu_40_in_2, msg_to_check_it_13_cnu_40_in_3, msg_to_check_it_13_cnu_40_in_4, msg_to_check_it_13_cnu_40_in_5, msg_to_check_it_13_cnu_41_in_0, msg_to_check_it_13_cnu_41_in_1, msg_to_check_it_13_cnu_41_in_2, msg_to_check_it_13_cnu_41_in_3, msg_to_check_it_13_cnu_41_in_4, msg_to_check_it_13_cnu_41_in_5, msg_to_check_it_13_cnu_42_in_0, msg_to_check_it_13_cnu_42_in_1, msg_to_check_it_13_cnu_42_in_2, msg_to_check_it_13_cnu_42_in_3, msg_to_check_it_13_cnu_42_in_4, msg_to_check_it_13_cnu_42_in_5, msg_to_check_it_13_cnu_43_in_0, msg_to_check_it_13_cnu_43_in_1, msg_to_check_it_13_cnu_43_in_2, msg_to_check_it_13_cnu_43_in_3, msg_to_check_it_13_cnu_43_in_4, msg_to_check_it_13_cnu_43_in_5, msg_to_check_it_13_cnu_44_in_0, msg_to_check_it_13_cnu_44_in_1, msg_to_check_it_13_cnu_44_in_2, msg_to_check_it_13_cnu_44_in_3, msg_to_check_it_13_cnu_44_in_4, msg_to_check_it_13_cnu_44_in_5, msg_to_check_it_13_cnu_45_in_0, msg_to_check_it_13_cnu_45_in_1, msg_to_check_it_13_cnu_45_in_2, msg_to_check_it_13_cnu_45_in_3, msg_to_check_it_13_cnu_45_in_4, msg_to_check_it_13_cnu_45_in_5, msg_to_check_it_13_cnu_46_in_0, msg_to_check_it_13_cnu_46_in_1, msg_to_check_it_13_cnu_46_in_2, msg_to_check_it_13_cnu_46_in_3, msg_to_check_it_13_cnu_46_in_4, msg_to_check_it_13_cnu_46_in_5, msg_to_check_it_13_cnu_47_in_0, msg_to_check_it_13_cnu_47_in_1, msg_to_check_it_13_cnu_47_in_2, msg_to_check_it_13_cnu_47_in_3, msg_to_check_it_13_cnu_47_in_4, msg_to_check_it_13_cnu_47_in_5, msg_to_check_it_13_cnu_48_in_0, msg_to_check_it_13_cnu_48_in_1, msg_to_check_it_13_cnu_48_in_2, msg_to_check_it_13_cnu_48_in_3, msg_to_check_it_13_cnu_48_in_4, msg_to_check_it_13_cnu_48_in_5, msg_to_check_it_13_cnu_49_in_0, msg_to_check_it_13_cnu_49_in_1, msg_to_check_it_13_cnu_49_in_2, msg_to_check_it_13_cnu_49_in_3, msg_to_check_it_13_cnu_49_in_4, msg_to_check_it_13_cnu_49_in_5, msg_to_check_it_13_cnu_50_in_0, msg_to_check_it_13_cnu_50_in_1, msg_to_check_it_13_cnu_50_in_2, msg_to_check_it_13_cnu_50_in_3, msg_to_check_it_13_cnu_50_in_4, msg_to_check_it_13_cnu_50_in_5, msg_to_check_it_13_cnu_51_in_0, msg_to_check_it_13_cnu_51_in_1, msg_to_check_it_13_cnu_51_in_2, msg_to_check_it_13_cnu_51_in_3, msg_to_check_it_13_cnu_51_in_4, msg_to_check_it_13_cnu_51_in_5, msg_to_check_it_13_cnu_52_in_0, msg_to_check_it_13_cnu_52_in_1, msg_to_check_it_13_cnu_52_in_2, msg_to_check_it_13_cnu_52_in_3, msg_to_check_it_13_cnu_52_in_4, msg_to_check_it_13_cnu_52_in_5, msg_to_check_it_13_cnu_53_in_0, msg_to_check_it_13_cnu_53_in_1, msg_to_check_it_13_cnu_53_in_2, msg_to_check_it_13_cnu_53_in_3, msg_to_check_it_13_cnu_53_in_4, msg_to_check_it_13_cnu_53_in_5, msg_to_check_it_13_cnu_54_in_0, msg_to_check_it_13_cnu_54_in_1, msg_to_check_it_13_cnu_54_in_2, msg_to_check_it_13_cnu_54_in_3, msg_to_check_it_13_cnu_54_in_4, msg_to_check_it_13_cnu_54_in_5, msg_to_check_it_13_cnu_55_in_0, msg_to_check_it_13_cnu_55_in_1, msg_to_check_it_13_cnu_55_in_2, msg_to_check_it_13_cnu_55_in_3, msg_to_check_it_13_cnu_55_in_4, msg_to_check_it_13_cnu_55_in_5, msg_to_check_it_13_cnu_56_in_0, msg_to_check_it_13_cnu_56_in_1, msg_to_check_it_13_cnu_56_in_2, msg_to_check_it_13_cnu_56_in_3, msg_to_check_it_13_cnu_56_in_4, msg_to_check_it_13_cnu_56_in_5, msg_to_check_it_13_cnu_57_in_0, msg_to_check_it_13_cnu_57_in_1, msg_to_check_it_13_cnu_57_in_2, msg_to_check_it_13_cnu_57_in_3, msg_to_check_it_13_cnu_57_in_4, msg_to_check_it_13_cnu_57_in_5, msg_to_check_it_13_cnu_58_in_0, msg_to_check_it_13_cnu_58_in_1, msg_to_check_it_13_cnu_58_in_2, msg_to_check_it_13_cnu_58_in_3, msg_to_check_it_13_cnu_58_in_4, msg_to_check_it_13_cnu_58_in_5, msg_to_check_it_13_cnu_59_in_0, msg_to_check_it_13_cnu_59_in_1, msg_to_check_it_13_cnu_59_in_2, msg_to_check_it_13_cnu_59_in_3, msg_to_check_it_13_cnu_59_in_4, msg_to_check_it_13_cnu_59_in_5, msg_to_check_it_13_cnu_60_in_0, msg_to_check_it_13_cnu_60_in_1, msg_to_check_it_13_cnu_60_in_2, msg_to_check_it_13_cnu_60_in_3, msg_to_check_it_13_cnu_60_in_4, msg_to_check_it_13_cnu_60_in_5, msg_to_check_it_13_cnu_61_in_0, msg_to_check_it_13_cnu_61_in_1, msg_to_check_it_13_cnu_61_in_2, msg_to_check_it_13_cnu_61_in_3, msg_to_check_it_13_cnu_61_in_4, msg_to_check_it_13_cnu_61_in_5, msg_to_check_it_13_cnu_62_in_0, msg_to_check_it_13_cnu_62_in_1, msg_to_check_it_13_cnu_62_in_2, msg_to_check_it_13_cnu_62_in_3, msg_to_check_it_13_cnu_62_in_4, msg_to_check_it_13_cnu_62_in_5, msg_to_check_it_13_cnu_63_in_0, msg_to_check_it_13_cnu_63_in_1, msg_to_check_it_13_cnu_63_in_2, msg_to_check_it_13_cnu_63_in_3, msg_to_check_it_13_cnu_63_in_4, msg_to_check_it_13_cnu_63_in_5, msg_to_check_it_13_cnu_64_in_0, msg_to_check_it_13_cnu_64_in_1, msg_to_check_it_13_cnu_64_in_2, msg_to_check_it_13_cnu_64_in_3, msg_to_check_it_13_cnu_64_in_4, msg_to_check_it_13_cnu_64_in_5, msg_to_check_it_13_cnu_65_in_0, msg_to_check_it_13_cnu_65_in_1, msg_to_check_it_13_cnu_65_in_2, msg_to_check_it_13_cnu_65_in_3, msg_to_check_it_13_cnu_65_in_4, msg_to_check_it_13_cnu_65_in_5, msg_to_check_it_13_cnu_66_in_0, msg_to_check_it_13_cnu_66_in_1, msg_to_check_it_13_cnu_66_in_2, msg_to_check_it_13_cnu_66_in_3, msg_to_check_it_13_cnu_66_in_4, msg_to_check_it_13_cnu_66_in_5, msg_to_check_it_13_cnu_67_in_0, msg_to_check_it_13_cnu_67_in_1, msg_to_check_it_13_cnu_67_in_2, msg_to_check_it_13_cnu_67_in_3, msg_to_check_it_13_cnu_67_in_4, msg_to_check_it_13_cnu_67_in_5, msg_to_check_it_13_cnu_68_in_0, msg_to_check_it_13_cnu_68_in_1, msg_to_check_it_13_cnu_68_in_2, msg_to_check_it_13_cnu_68_in_3, msg_to_check_it_13_cnu_68_in_4, msg_to_check_it_13_cnu_68_in_5, msg_to_check_it_13_cnu_69_in_0, msg_to_check_it_13_cnu_69_in_1, msg_to_check_it_13_cnu_69_in_2, msg_to_check_it_13_cnu_69_in_3, msg_to_check_it_13_cnu_69_in_4, msg_to_check_it_13_cnu_69_in_5, msg_to_check_it_13_cnu_70_in_0, msg_to_check_it_13_cnu_70_in_1, msg_to_check_it_13_cnu_70_in_2, msg_to_check_it_13_cnu_70_in_3, msg_to_check_it_13_cnu_70_in_4, msg_to_check_it_13_cnu_70_in_5, msg_to_check_it_13_cnu_71_in_0, msg_to_check_it_13_cnu_71_in_1, msg_to_check_it_13_cnu_71_in_2, msg_to_check_it_13_cnu_71_in_3, msg_to_check_it_13_cnu_71_in_4, msg_to_check_it_13_cnu_71_in_5, msg_to_check_it_13_cnu_72_in_0, msg_to_check_it_13_cnu_72_in_1, msg_to_check_it_13_cnu_72_in_2, msg_to_check_it_13_cnu_72_in_3, msg_to_check_it_13_cnu_72_in_4, msg_to_check_it_13_cnu_72_in_5, msg_to_check_it_13_cnu_73_in_0, msg_to_check_it_13_cnu_73_in_1, msg_to_check_it_13_cnu_73_in_2, msg_to_check_it_13_cnu_73_in_3, msg_to_check_it_13_cnu_73_in_4, msg_to_check_it_13_cnu_73_in_5, msg_to_check_it_13_cnu_74_in_0, msg_to_check_it_13_cnu_74_in_1, msg_to_check_it_13_cnu_74_in_2, msg_to_check_it_13_cnu_74_in_3, msg_to_check_it_13_cnu_74_in_4, msg_to_check_it_13_cnu_74_in_5, msg_to_check_it_13_cnu_75_in_0, msg_to_check_it_13_cnu_75_in_1, msg_to_check_it_13_cnu_75_in_2, msg_to_check_it_13_cnu_75_in_3, msg_to_check_it_13_cnu_75_in_4, msg_to_check_it_13_cnu_75_in_5, msg_to_check_it_13_cnu_76_in_0, msg_to_check_it_13_cnu_76_in_1, msg_to_check_it_13_cnu_76_in_2, msg_to_check_it_13_cnu_76_in_3, msg_to_check_it_13_cnu_76_in_4, msg_to_check_it_13_cnu_76_in_5, msg_to_check_it_13_cnu_77_in_0, msg_to_check_it_13_cnu_77_in_1, msg_to_check_it_13_cnu_77_in_2, msg_to_check_it_13_cnu_77_in_3, msg_to_check_it_13_cnu_77_in_4, msg_to_check_it_13_cnu_77_in_5, msg_to_check_it_13_cnu_78_in_0, msg_to_check_it_13_cnu_78_in_1, msg_to_check_it_13_cnu_78_in_2, msg_to_check_it_13_cnu_78_in_3, msg_to_check_it_13_cnu_78_in_4, msg_to_check_it_13_cnu_78_in_5, msg_to_check_it_13_cnu_79_in_0, msg_to_check_it_13_cnu_79_in_1, msg_to_check_it_13_cnu_79_in_2, msg_to_check_it_13_cnu_79_in_3, msg_to_check_it_13_cnu_79_in_4, msg_to_check_it_13_cnu_79_in_5, msg_to_check_it_13_cnu_80_in_0, msg_to_check_it_13_cnu_80_in_1, msg_to_check_it_13_cnu_80_in_2, msg_to_check_it_13_cnu_80_in_3, msg_to_check_it_13_cnu_80_in_4, msg_to_check_it_13_cnu_80_in_5, msg_to_check_it_13_cnu_81_in_0, msg_to_check_it_13_cnu_81_in_1, msg_to_check_it_13_cnu_81_in_2, msg_to_check_it_13_cnu_81_in_3, msg_to_check_it_13_cnu_81_in_4, msg_to_check_it_13_cnu_81_in_5, msg_to_check_it_13_cnu_82_in_0, msg_to_check_it_13_cnu_82_in_1, msg_to_check_it_13_cnu_82_in_2, msg_to_check_it_13_cnu_82_in_3, msg_to_check_it_13_cnu_82_in_4, msg_to_check_it_13_cnu_82_in_5, msg_to_check_it_13_cnu_83_in_0, msg_to_check_it_13_cnu_83_in_1, msg_to_check_it_13_cnu_83_in_2, msg_to_check_it_13_cnu_83_in_3, msg_to_check_it_13_cnu_83_in_4, msg_to_check_it_13_cnu_83_in_5, msg_to_check_it_13_cnu_84_in_0, msg_to_check_it_13_cnu_84_in_1, msg_to_check_it_13_cnu_84_in_2, msg_to_check_it_13_cnu_84_in_3, msg_to_check_it_13_cnu_84_in_4, msg_to_check_it_13_cnu_84_in_5, msg_to_check_it_13_cnu_85_in_0, msg_to_check_it_13_cnu_85_in_1, msg_to_check_it_13_cnu_85_in_2, msg_to_check_it_13_cnu_85_in_3, msg_to_check_it_13_cnu_85_in_4, msg_to_check_it_13_cnu_85_in_5, msg_to_check_it_13_cnu_86_in_0, msg_to_check_it_13_cnu_86_in_1, msg_to_check_it_13_cnu_86_in_2, msg_to_check_it_13_cnu_86_in_3, msg_to_check_it_13_cnu_86_in_4, msg_to_check_it_13_cnu_86_in_5, msg_to_check_it_13_cnu_87_in_0, msg_to_check_it_13_cnu_87_in_1, msg_to_check_it_13_cnu_87_in_2, msg_to_check_it_13_cnu_87_in_3, msg_to_check_it_13_cnu_87_in_4, msg_to_check_it_13_cnu_87_in_5, msg_to_check_it_13_cnu_88_in_0, msg_to_check_it_13_cnu_88_in_1, msg_to_check_it_13_cnu_88_in_2, msg_to_check_it_13_cnu_88_in_3, msg_to_check_it_13_cnu_88_in_4, msg_to_check_it_13_cnu_88_in_5, msg_to_check_it_13_cnu_89_in_0, msg_to_check_it_13_cnu_89_in_1, msg_to_check_it_13_cnu_89_in_2, msg_to_check_it_13_cnu_89_in_3, msg_to_check_it_13_cnu_89_in_4, msg_to_check_it_13_cnu_89_in_5, msg_to_check_it_13_cnu_90_in_0, msg_to_check_it_13_cnu_90_in_1, msg_to_check_it_13_cnu_90_in_2, msg_to_check_it_13_cnu_90_in_3, msg_to_check_it_13_cnu_90_in_4, msg_to_check_it_13_cnu_90_in_5, msg_to_check_it_13_cnu_91_in_0, msg_to_check_it_13_cnu_91_in_1, msg_to_check_it_13_cnu_91_in_2, msg_to_check_it_13_cnu_91_in_3, msg_to_check_it_13_cnu_91_in_4, msg_to_check_it_13_cnu_91_in_5, msg_to_check_it_13_cnu_92_in_0, msg_to_check_it_13_cnu_92_in_1, msg_to_check_it_13_cnu_92_in_2, msg_to_check_it_13_cnu_92_in_3, msg_to_check_it_13_cnu_92_in_4, msg_to_check_it_13_cnu_92_in_5, msg_to_check_it_13_cnu_93_in_0, msg_to_check_it_13_cnu_93_in_1, msg_to_check_it_13_cnu_93_in_2, msg_to_check_it_13_cnu_93_in_3, msg_to_check_it_13_cnu_93_in_4, msg_to_check_it_13_cnu_93_in_5, msg_to_check_it_13_cnu_94_in_0, msg_to_check_it_13_cnu_94_in_1, msg_to_check_it_13_cnu_94_in_2, msg_to_check_it_13_cnu_94_in_3, msg_to_check_it_13_cnu_94_in_4, msg_to_check_it_13_cnu_94_in_5, msg_to_check_it_13_cnu_95_in_0, msg_to_check_it_13_cnu_95_in_1, msg_to_check_it_13_cnu_95_in_2, msg_to_check_it_13_cnu_95_in_3, msg_to_check_it_13_cnu_95_in_4, msg_to_check_it_13_cnu_95_in_5, msg_to_check_it_13_cnu_96_in_0, msg_to_check_it_13_cnu_96_in_1, msg_to_check_it_13_cnu_96_in_2, msg_to_check_it_13_cnu_96_in_3, msg_to_check_it_13_cnu_96_in_4, msg_to_check_it_13_cnu_96_in_5, msg_to_check_it_13_cnu_97_in_0, msg_to_check_it_13_cnu_97_in_1, msg_to_check_it_13_cnu_97_in_2, msg_to_check_it_13_cnu_97_in_3, msg_to_check_it_13_cnu_97_in_4, msg_to_check_it_13_cnu_97_in_5, msg_to_check_it_13_cnu_98_in_0, msg_to_check_it_13_cnu_98_in_1, msg_to_check_it_13_cnu_98_in_2, msg_to_check_it_13_cnu_98_in_3, msg_to_check_it_13_cnu_98_in_4, msg_to_check_it_13_cnu_98_in_5, msg_to_check_it_14_cnu_0_in_0, msg_to_check_it_14_cnu_0_in_1, msg_to_check_it_14_cnu_0_in_2, msg_to_check_it_14_cnu_0_in_3, msg_to_check_it_14_cnu_0_in_4, msg_to_check_it_14_cnu_0_in_5, msg_to_check_it_14_cnu_1_in_0, msg_to_check_it_14_cnu_1_in_1, msg_to_check_it_14_cnu_1_in_2, msg_to_check_it_14_cnu_1_in_3, msg_to_check_it_14_cnu_1_in_4, msg_to_check_it_14_cnu_1_in_5, msg_to_check_it_14_cnu_2_in_0, msg_to_check_it_14_cnu_2_in_1, msg_to_check_it_14_cnu_2_in_2, msg_to_check_it_14_cnu_2_in_3, msg_to_check_it_14_cnu_2_in_4, msg_to_check_it_14_cnu_2_in_5, msg_to_check_it_14_cnu_3_in_0, msg_to_check_it_14_cnu_3_in_1, msg_to_check_it_14_cnu_3_in_2, msg_to_check_it_14_cnu_3_in_3, msg_to_check_it_14_cnu_3_in_4, msg_to_check_it_14_cnu_3_in_5, msg_to_check_it_14_cnu_4_in_0, msg_to_check_it_14_cnu_4_in_1, msg_to_check_it_14_cnu_4_in_2, msg_to_check_it_14_cnu_4_in_3, msg_to_check_it_14_cnu_4_in_4, msg_to_check_it_14_cnu_4_in_5, msg_to_check_it_14_cnu_5_in_0, msg_to_check_it_14_cnu_5_in_1, msg_to_check_it_14_cnu_5_in_2, msg_to_check_it_14_cnu_5_in_3, msg_to_check_it_14_cnu_5_in_4, msg_to_check_it_14_cnu_5_in_5, msg_to_check_it_14_cnu_6_in_0, msg_to_check_it_14_cnu_6_in_1, msg_to_check_it_14_cnu_6_in_2, msg_to_check_it_14_cnu_6_in_3, msg_to_check_it_14_cnu_6_in_4, msg_to_check_it_14_cnu_6_in_5, msg_to_check_it_14_cnu_7_in_0, msg_to_check_it_14_cnu_7_in_1, msg_to_check_it_14_cnu_7_in_2, msg_to_check_it_14_cnu_7_in_3, msg_to_check_it_14_cnu_7_in_4, msg_to_check_it_14_cnu_7_in_5, msg_to_check_it_14_cnu_8_in_0, msg_to_check_it_14_cnu_8_in_1, msg_to_check_it_14_cnu_8_in_2, msg_to_check_it_14_cnu_8_in_3, msg_to_check_it_14_cnu_8_in_4, msg_to_check_it_14_cnu_8_in_5, msg_to_check_it_14_cnu_9_in_0, msg_to_check_it_14_cnu_9_in_1, msg_to_check_it_14_cnu_9_in_2, msg_to_check_it_14_cnu_9_in_3, msg_to_check_it_14_cnu_9_in_4, msg_to_check_it_14_cnu_9_in_5, msg_to_check_it_14_cnu_10_in_0, msg_to_check_it_14_cnu_10_in_1, msg_to_check_it_14_cnu_10_in_2, msg_to_check_it_14_cnu_10_in_3, msg_to_check_it_14_cnu_10_in_4, msg_to_check_it_14_cnu_10_in_5, msg_to_check_it_14_cnu_11_in_0, msg_to_check_it_14_cnu_11_in_1, msg_to_check_it_14_cnu_11_in_2, msg_to_check_it_14_cnu_11_in_3, msg_to_check_it_14_cnu_11_in_4, msg_to_check_it_14_cnu_11_in_5, msg_to_check_it_14_cnu_12_in_0, msg_to_check_it_14_cnu_12_in_1, msg_to_check_it_14_cnu_12_in_2, msg_to_check_it_14_cnu_12_in_3, msg_to_check_it_14_cnu_12_in_4, msg_to_check_it_14_cnu_12_in_5, msg_to_check_it_14_cnu_13_in_0, msg_to_check_it_14_cnu_13_in_1, msg_to_check_it_14_cnu_13_in_2, msg_to_check_it_14_cnu_13_in_3, msg_to_check_it_14_cnu_13_in_4, msg_to_check_it_14_cnu_13_in_5, msg_to_check_it_14_cnu_14_in_0, msg_to_check_it_14_cnu_14_in_1, msg_to_check_it_14_cnu_14_in_2, msg_to_check_it_14_cnu_14_in_3, msg_to_check_it_14_cnu_14_in_4, msg_to_check_it_14_cnu_14_in_5, msg_to_check_it_14_cnu_15_in_0, msg_to_check_it_14_cnu_15_in_1, msg_to_check_it_14_cnu_15_in_2, msg_to_check_it_14_cnu_15_in_3, msg_to_check_it_14_cnu_15_in_4, msg_to_check_it_14_cnu_15_in_5, msg_to_check_it_14_cnu_16_in_0, msg_to_check_it_14_cnu_16_in_1, msg_to_check_it_14_cnu_16_in_2, msg_to_check_it_14_cnu_16_in_3, msg_to_check_it_14_cnu_16_in_4, msg_to_check_it_14_cnu_16_in_5, msg_to_check_it_14_cnu_17_in_0, msg_to_check_it_14_cnu_17_in_1, msg_to_check_it_14_cnu_17_in_2, msg_to_check_it_14_cnu_17_in_3, msg_to_check_it_14_cnu_17_in_4, msg_to_check_it_14_cnu_17_in_5, msg_to_check_it_14_cnu_18_in_0, msg_to_check_it_14_cnu_18_in_1, msg_to_check_it_14_cnu_18_in_2, msg_to_check_it_14_cnu_18_in_3, msg_to_check_it_14_cnu_18_in_4, msg_to_check_it_14_cnu_18_in_5, msg_to_check_it_14_cnu_19_in_0, msg_to_check_it_14_cnu_19_in_1, msg_to_check_it_14_cnu_19_in_2, msg_to_check_it_14_cnu_19_in_3, msg_to_check_it_14_cnu_19_in_4, msg_to_check_it_14_cnu_19_in_5, msg_to_check_it_14_cnu_20_in_0, msg_to_check_it_14_cnu_20_in_1, msg_to_check_it_14_cnu_20_in_2, msg_to_check_it_14_cnu_20_in_3, msg_to_check_it_14_cnu_20_in_4, msg_to_check_it_14_cnu_20_in_5, msg_to_check_it_14_cnu_21_in_0, msg_to_check_it_14_cnu_21_in_1, msg_to_check_it_14_cnu_21_in_2, msg_to_check_it_14_cnu_21_in_3, msg_to_check_it_14_cnu_21_in_4, msg_to_check_it_14_cnu_21_in_5, msg_to_check_it_14_cnu_22_in_0, msg_to_check_it_14_cnu_22_in_1, msg_to_check_it_14_cnu_22_in_2, msg_to_check_it_14_cnu_22_in_3, msg_to_check_it_14_cnu_22_in_4, msg_to_check_it_14_cnu_22_in_5, msg_to_check_it_14_cnu_23_in_0, msg_to_check_it_14_cnu_23_in_1, msg_to_check_it_14_cnu_23_in_2, msg_to_check_it_14_cnu_23_in_3, msg_to_check_it_14_cnu_23_in_4, msg_to_check_it_14_cnu_23_in_5, msg_to_check_it_14_cnu_24_in_0, msg_to_check_it_14_cnu_24_in_1, msg_to_check_it_14_cnu_24_in_2, msg_to_check_it_14_cnu_24_in_3, msg_to_check_it_14_cnu_24_in_4, msg_to_check_it_14_cnu_24_in_5, msg_to_check_it_14_cnu_25_in_0, msg_to_check_it_14_cnu_25_in_1, msg_to_check_it_14_cnu_25_in_2, msg_to_check_it_14_cnu_25_in_3, msg_to_check_it_14_cnu_25_in_4, msg_to_check_it_14_cnu_25_in_5, msg_to_check_it_14_cnu_26_in_0, msg_to_check_it_14_cnu_26_in_1, msg_to_check_it_14_cnu_26_in_2, msg_to_check_it_14_cnu_26_in_3, msg_to_check_it_14_cnu_26_in_4, msg_to_check_it_14_cnu_26_in_5, msg_to_check_it_14_cnu_27_in_0, msg_to_check_it_14_cnu_27_in_1, msg_to_check_it_14_cnu_27_in_2, msg_to_check_it_14_cnu_27_in_3, msg_to_check_it_14_cnu_27_in_4, msg_to_check_it_14_cnu_27_in_5, msg_to_check_it_14_cnu_28_in_0, msg_to_check_it_14_cnu_28_in_1, msg_to_check_it_14_cnu_28_in_2, msg_to_check_it_14_cnu_28_in_3, msg_to_check_it_14_cnu_28_in_4, msg_to_check_it_14_cnu_28_in_5, msg_to_check_it_14_cnu_29_in_0, msg_to_check_it_14_cnu_29_in_1, msg_to_check_it_14_cnu_29_in_2, msg_to_check_it_14_cnu_29_in_3, msg_to_check_it_14_cnu_29_in_4, msg_to_check_it_14_cnu_29_in_5, msg_to_check_it_14_cnu_30_in_0, msg_to_check_it_14_cnu_30_in_1, msg_to_check_it_14_cnu_30_in_2, msg_to_check_it_14_cnu_30_in_3, msg_to_check_it_14_cnu_30_in_4, msg_to_check_it_14_cnu_30_in_5, msg_to_check_it_14_cnu_31_in_0, msg_to_check_it_14_cnu_31_in_1, msg_to_check_it_14_cnu_31_in_2, msg_to_check_it_14_cnu_31_in_3, msg_to_check_it_14_cnu_31_in_4, msg_to_check_it_14_cnu_31_in_5, msg_to_check_it_14_cnu_32_in_0, msg_to_check_it_14_cnu_32_in_1, msg_to_check_it_14_cnu_32_in_2, msg_to_check_it_14_cnu_32_in_3, msg_to_check_it_14_cnu_32_in_4, msg_to_check_it_14_cnu_32_in_5, msg_to_check_it_14_cnu_33_in_0, msg_to_check_it_14_cnu_33_in_1, msg_to_check_it_14_cnu_33_in_2, msg_to_check_it_14_cnu_33_in_3, msg_to_check_it_14_cnu_33_in_4, msg_to_check_it_14_cnu_33_in_5, msg_to_check_it_14_cnu_34_in_0, msg_to_check_it_14_cnu_34_in_1, msg_to_check_it_14_cnu_34_in_2, msg_to_check_it_14_cnu_34_in_3, msg_to_check_it_14_cnu_34_in_4, msg_to_check_it_14_cnu_34_in_5, msg_to_check_it_14_cnu_35_in_0, msg_to_check_it_14_cnu_35_in_1, msg_to_check_it_14_cnu_35_in_2, msg_to_check_it_14_cnu_35_in_3, msg_to_check_it_14_cnu_35_in_4, msg_to_check_it_14_cnu_35_in_5, msg_to_check_it_14_cnu_36_in_0, msg_to_check_it_14_cnu_36_in_1, msg_to_check_it_14_cnu_36_in_2, msg_to_check_it_14_cnu_36_in_3, msg_to_check_it_14_cnu_36_in_4, msg_to_check_it_14_cnu_36_in_5, msg_to_check_it_14_cnu_37_in_0, msg_to_check_it_14_cnu_37_in_1, msg_to_check_it_14_cnu_37_in_2, msg_to_check_it_14_cnu_37_in_3, msg_to_check_it_14_cnu_37_in_4, msg_to_check_it_14_cnu_37_in_5, msg_to_check_it_14_cnu_38_in_0, msg_to_check_it_14_cnu_38_in_1, msg_to_check_it_14_cnu_38_in_2, msg_to_check_it_14_cnu_38_in_3, msg_to_check_it_14_cnu_38_in_4, msg_to_check_it_14_cnu_38_in_5, msg_to_check_it_14_cnu_39_in_0, msg_to_check_it_14_cnu_39_in_1, msg_to_check_it_14_cnu_39_in_2, msg_to_check_it_14_cnu_39_in_3, msg_to_check_it_14_cnu_39_in_4, msg_to_check_it_14_cnu_39_in_5, msg_to_check_it_14_cnu_40_in_0, msg_to_check_it_14_cnu_40_in_1, msg_to_check_it_14_cnu_40_in_2, msg_to_check_it_14_cnu_40_in_3, msg_to_check_it_14_cnu_40_in_4, msg_to_check_it_14_cnu_40_in_5, msg_to_check_it_14_cnu_41_in_0, msg_to_check_it_14_cnu_41_in_1, msg_to_check_it_14_cnu_41_in_2, msg_to_check_it_14_cnu_41_in_3, msg_to_check_it_14_cnu_41_in_4, msg_to_check_it_14_cnu_41_in_5, msg_to_check_it_14_cnu_42_in_0, msg_to_check_it_14_cnu_42_in_1, msg_to_check_it_14_cnu_42_in_2, msg_to_check_it_14_cnu_42_in_3, msg_to_check_it_14_cnu_42_in_4, msg_to_check_it_14_cnu_42_in_5, msg_to_check_it_14_cnu_43_in_0, msg_to_check_it_14_cnu_43_in_1, msg_to_check_it_14_cnu_43_in_2, msg_to_check_it_14_cnu_43_in_3, msg_to_check_it_14_cnu_43_in_4, msg_to_check_it_14_cnu_43_in_5, msg_to_check_it_14_cnu_44_in_0, msg_to_check_it_14_cnu_44_in_1, msg_to_check_it_14_cnu_44_in_2, msg_to_check_it_14_cnu_44_in_3, msg_to_check_it_14_cnu_44_in_4, msg_to_check_it_14_cnu_44_in_5, msg_to_check_it_14_cnu_45_in_0, msg_to_check_it_14_cnu_45_in_1, msg_to_check_it_14_cnu_45_in_2, msg_to_check_it_14_cnu_45_in_3, msg_to_check_it_14_cnu_45_in_4, msg_to_check_it_14_cnu_45_in_5, msg_to_check_it_14_cnu_46_in_0, msg_to_check_it_14_cnu_46_in_1, msg_to_check_it_14_cnu_46_in_2, msg_to_check_it_14_cnu_46_in_3, msg_to_check_it_14_cnu_46_in_4, msg_to_check_it_14_cnu_46_in_5, msg_to_check_it_14_cnu_47_in_0, msg_to_check_it_14_cnu_47_in_1, msg_to_check_it_14_cnu_47_in_2, msg_to_check_it_14_cnu_47_in_3, msg_to_check_it_14_cnu_47_in_4, msg_to_check_it_14_cnu_47_in_5, msg_to_check_it_14_cnu_48_in_0, msg_to_check_it_14_cnu_48_in_1, msg_to_check_it_14_cnu_48_in_2, msg_to_check_it_14_cnu_48_in_3, msg_to_check_it_14_cnu_48_in_4, msg_to_check_it_14_cnu_48_in_5, msg_to_check_it_14_cnu_49_in_0, msg_to_check_it_14_cnu_49_in_1, msg_to_check_it_14_cnu_49_in_2, msg_to_check_it_14_cnu_49_in_3, msg_to_check_it_14_cnu_49_in_4, msg_to_check_it_14_cnu_49_in_5, msg_to_check_it_14_cnu_50_in_0, msg_to_check_it_14_cnu_50_in_1, msg_to_check_it_14_cnu_50_in_2, msg_to_check_it_14_cnu_50_in_3, msg_to_check_it_14_cnu_50_in_4, msg_to_check_it_14_cnu_50_in_5, msg_to_check_it_14_cnu_51_in_0, msg_to_check_it_14_cnu_51_in_1, msg_to_check_it_14_cnu_51_in_2, msg_to_check_it_14_cnu_51_in_3, msg_to_check_it_14_cnu_51_in_4, msg_to_check_it_14_cnu_51_in_5, msg_to_check_it_14_cnu_52_in_0, msg_to_check_it_14_cnu_52_in_1, msg_to_check_it_14_cnu_52_in_2, msg_to_check_it_14_cnu_52_in_3, msg_to_check_it_14_cnu_52_in_4, msg_to_check_it_14_cnu_52_in_5, msg_to_check_it_14_cnu_53_in_0, msg_to_check_it_14_cnu_53_in_1, msg_to_check_it_14_cnu_53_in_2, msg_to_check_it_14_cnu_53_in_3, msg_to_check_it_14_cnu_53_in_4, msg_to_check_it_14_cnu_53_in_5, msg_to_check_it_14_cnu_54_in_0, msg_to_check_it_14_cnu_54_in_1, msg_to_check_it_14_cnu_54_in_2, msg_to_check_it_14_cnu_54_in_3, msg_to_check_it_14_cnu_54_in_4, msg_to_check_it_14_cnu_54_in_5, msg_to_check_it_14_cnu_55_in_0, msg_to_check_it_14_cnu_55_in_1, msg_to_check_it_14_cnu_55_in_2, msg_to_check_it_14_cnu_55_in_3, msg_to_check_it_14_cnu_55_in_4, msg_to_check_it_14_cnu_55_in_5, msg_to_check_it_14_cnu_56_in_0, msg_to_check_it_14_cnu_56_in_1, msg_to_check_it_14_cnu_56_in_2, msg_to_check_it_14_cnu_56_in_3, msg_to_check_it_14_cnu_56_in_4, msg_to_check_it_14_cnu_56_in_5, msg_to_check_it_14_cnu_57_in_0, msg_to_check_it_14_cnu_57_in_1, msg_to_check_it_14_cnu_57_in_2, msg_to_check_it_14_cnu_57_in_3, msg_to_check_it_14_cnu_57_in_4, msg_to_check_it_14_cnu_57_in_5, msg_to_check_it_14_cnu_58_in_0, msg_to_check_it_14_cnu_58_in_1, msg_to_check_it_14_cnu_58_in_2, msg_to_check_it_14_cnu_58_in_3, msg_to_check_it_14_cnu_58_in_4, msg_to_check_it_14_cnu_58_in_5, msg_to_check_it_14_cnu_59_in_0, msg_to_check_it_14_cnu_59_in_1, msg_to_check_it_14_cnu_59_in_2, msg_to_check_it_14_cnu_59_in_3, msg_to_check_it_14_cnu_59_in_4, msg_to_check_it_14_cnu_59_in_5, msg_to_check_it_14_cnu_60_in_0, msg_to_check_it_14_cnu_60_in_1, msg_to_check_it_14_cnu_60_in_2, msg_to_check_it_14_cnu_60_in_3, msg_to_check_it_14_cnu_60_in_4, msg_to_check_it_14_cnu_60_in_5, msg_to_check_it_14_cnu_61_in_0, msg_to_check_it_14_cnu_61_in_1, msg_to_check_it_14_cnu_61_in_2, msg_to_check_it_14_cnu_61_in_3, msg_to_check_it_14_cnu_61_in_4, msg_to_check_it_14_cnu_61_in_5, msg_to_check_it_14_cnu_62_in_0, msg_to_check_it_14_cnu_62_in_1, msg_to_check_it_14_cnu_62_in_2, msg_to_check_it_14_cnu_62_in_3, msg_to_check_it_14_cnu_62_in_4, msg_to_check_it_14_cnu_62_in_5, msg_to_check_it_14_cnu_63_in_0, msg_to_check_it_14_cnu_63_in_1, msg_to_check_it_14_cnu_63_in_2, msg_to_check_it_14_cnu_63_in_3, msg_to_check_it_14_cnu_63_in_4, msg_to_check_it_14_cnu_63_in_5, msg_to_check_it_14_cnu_64_in_0, msg_to_check_it_14_cnu_64_in_1, msg_to_check_it_14_cnu_64_in_2, msg_to_check_it_14_cnu_64_in_3, msg_to_check_it_14_cnu_64_in_4, msg_to_check_it_14_cnu_64_in_5, msg_to_check_it_14_cnu_65_in_0, msg_to_check_it_14_cnu_65_in_1, msg_to_check_it_14_cnu_65_in_2, msg_to_check_it_14_cnu_65_in_3, msg_to_check_it_14_cnu_65_in_4, msg_to_check_it_14_cnu_65_in_5, msg_to_check_it_14_cnu_66_in_0, msg_to_check_it_14_cnu_66_in_1, msg_to_check_it_14_cnu_66_in_2, msg_to_check_it_14_cnu_66_in_3, msg_to_check_it_14_cnu_66_in_4, msg_to_check_it_14_cnu_66_in_5, msg_to_check_it_14_cnu_67_in_0, msg_to_check_it_14_cnu_67_in_1, msg_to_check_it_14_cnu_67_in_2, msg_to_check_it_14_cnu_67_in_3, msg_to_check_it_14_cnu_67_in_4, msg_to_check_it_14_cnu_67_in_5, msg_to_check_it_14_cnu_68_in_0, msg_to_check_it_14_cnu_68_in_1, msg_to_check_it_14_cnu_68_in_2, msg_to_check_it_14_cnu_68_in_3, msg_to_check_it_14_cnu_68_in_4, msg_to_check_it_14_cnu_68_in_5, msg_to_check_it_14_cnu_69_in_0, msg_to_check_it_14_cnu_69_in_1, msg_to_check_it_14_cnu_69_in_2, msg_to_check_it_14_cnu_69_in_3, msg_to_check_it_14_cnu_69_in_4, msg_to_check_it_14_cnu_69_in_5, msg_to_check_it_14_cnu_70_in_0, msg_to_check_it_14_cnu_70_in_1, msg_to_check_it_14_cnu_70_in_2, msg_to_check_it_14_cnu_70_in_3, msg_to_check_it_14_cnu_70_in_4, msg_to_check_it_14_cnu_70_in_5, msg_to_check_it_14_cnu_71_in_0, msg_to_check_it_14_cnu_71_in_1, msg_to_check_it_14_cnu_71_in_2, msg_to_check_it_14_cnu_71_in_3, msg_to_check_it_14_cnu_71_in_4, msg_to_check_it_14_cnu_71_in_5, msg_to_check_it_14_cnu_72_in_0, msg_to_check_it_14_cnu_72_in_1, msg_to_check_it_14_cnu_72_in_2, msg_to_check_it_14_cnu_72_in_3, msg_to_check_it_14_cnu_72_in_4, msg_to_check_it_14_cnu_72_in_5, msg_to_check_it_14_cnu_73_in_0, msg_to_check_it_14_cnu_73_in_1, msg_to_check_it_14_cnu_73_in_2, msg_to_check_it_14_cnu_73_in_3, msg_to_check_it_14_cnu_73_in_4, msg_to_check_it_14_cnu_73_in_5, msg_to_check_it_14_cnu_74_in_0, msg_to_check_it_14_cnu_74_in_1, msg_to_check_it_14_cnu_74_in_2, msg_to_check_it_14_cnu_74_in_3, msg_to_check_it_14_cnu_74_in_4, msg_to_check_it_14_cnu_74_in_5, msg_to_check_it_14_cnu_75_in_0, msg_to_check_it_14_cnu_75_in_1, msg_to_check_it_14_cnu_75_in_2, msg_to_check_it_14_cnu_75_in_3, msg_to_check_it_14_cnu_75_in_4, msg_to_check_it_14_cnu_75_in_5, msg_to_check_it_14_cnu_76_in_0, msg_to_check_it_14_cnu_76_in_1, msg_to_check_it_14_cnu_76_in_2, msg_to_check_it_14_cnu_76_in_3, msg_to_check_it_14_cnu_76_in_4, msg_to_check_it_14_cnu_76_in_5, msg_to_check_it_14_cnu_77_in_0, msg_to_check_it_14_cnu_77_in_1, msg_to_check_it_14_cnu_77_in_2, msg_to_check_it_14_cnu_77_in_3, msg_to_check_it_14_cnu_77_in_4, msg_to_check_it_14_cnu_77_in_5, msg_to_check_it_14_cnu_78_in_0, msg_to_check_it_14_cnu_78_in_1, msg_to_check_it_14_cnu_78_in_2, msg_to_check_it_14_cnu_78_in_3, msg_to_check_it_14_cnu_78_in_4, msg_to_check_it_14_cnu_78_in_5, msg_to_check_it_14_cnu_79_in_0, msg_to_check_it_14_cnu_79_in_1, msg_to_check_it_14_cnu_79_in_2, msg_to_check_it_14_cnu_79_in_3, msg_to_check_it_14_cnu_79_in_4, msg_to_check_it_14_cnu_79_in_5, msg_to_check_it_14_cnu_80_in_0, msg_to_check_it_14_cnu_80_in_1, msg_to_check_it_14_cnu_80_in_2, msg_to_check_it_14_cnu_80_in_3, msg_to_check_it_14_cnu_80_in_4, msg_to_check_it_14_cnu_80_in_5, msg_to_check_it_14_cnu_81_in_0, msg_to_check_it_14_cnu_81_in_1, msg_to_check_it_14_cnu_81_in_2, msg_to_check_it_14_cnu_81_in_3, msg_to_check_it_14_cnu_81_in_4, msg_to_check_it_14_cnu_81_in_5, msg_to_check_it_14_cnu_82_in_0, msg_to_check_it_14_cnu_82_in_1, msg_to_check_it_14_cnu_82_in_2, msg_to_check_it_14_cnu_82_in_3, msg_to_check_it_14_cnu_82_in_4, msg_to_check_it_14_cnu_82_in_5, msg_to_check_it_14_cnu_83_in_0, msg_to_check_it_14_cnu_83_in_1, msg_to_check_it_14_cnu_83_in_2, msg_to_check_it_14_cnu_83_in_3, msg_to_check_it_14_cnu_83_in_4, msg_to_check_it_14_cnu_83_in_5, msg_to_check_it_14_cnu_84_in_0, msg_to_check_it_14_cnu_84_in_1, msg_to_check_it_14_cnu_84_in_2, msg_to_check_it_14_cnu_84_in_3, msg_to_check_it_14_cnu_84_in_4, msg_to_check_it_14_cnu_84_in_5, msg_to_check_it_14_cnu_85_in_0, msg_to_check_it_14_cnu_85_in_1, msg_to_check_it_14_cnu_85_in_2, msg_to_check_it_14_cnu_85_in_3, msg_to_check_it_14_cnu_85_in_4, msg_to_check_it_14_cnu_85_in_5, msg_to_check_it_14_cnu_86_in_0, msg_to_check_it_14_cnu_86_in_1, msg_to_check_it_14_cnu_86_in_2, msg_to_check_it_14_cnu_86_in_3, msg_to_check_it_14_cnu_86_in_4, msg_to_check_it_14_cnu_86_in_5, msg_to_check_it_14_cnu_87_in_0, msg_to_check_it_14_cnu_87_in_1, msg_to_check_it_14_cnu_87_in_2, msg_to_check_it_14_cnu_87_in_3, msg_to_check_it_14_cnu_87_in_4, msg_to_check_it_14_cnu_87_in_5, msg_to_check_it_14_cnu_88_in_0, msg_to_check_it_14_cnu_88_in_1, msg_to_check_it_14_cnu_88_in_2, msg_to_check_it_14_cnu_88_in_3, msg_to_check_it_14_cnu_88_in_4, msg_to_check_it_14_cnu_88_in_5, msg_to_check_it_14_cnu_89_in_0, msg_to_check_it_14_cnu_89_in_1, msg_to_check_it_14_cnu_89_in_2, msg_to_check_it_14_cnu_89_in_3, msg_to_check_it_14_cnu_89_in_4, msg_to_check_it_14_cnu_89_in_5, msg_to_check_it_14_cnu_90_in_0, msg_to_check_it_14_cnu_90_in_1, msg_to_check_it_14_cnu_90_in_2, msg_to_check_it_14_cnu_90_in_3, msg_to_check_it_14_cnu_90_in_4, msg_to_check_it_14_cnu_90_in_5, msg_to_check_it_14_cnu_91_in_0, msg_to_check_it_14_cnu_91_in_1, msg_to_check_it_14_cnu_91_in_2, msg_to_check_it_14_cnu_91_in_3, msg_to_check_it_14_cnu_91_in_4, msg_to_check_it_14_cnu_91_in_5, msg_to_check_it_14_cnu_92_in_0, msg_to_check_it_14_cnu_92_in_1, msg_to_check_it_14_cnu_92_in_2, msg_to_check_it_14_cnu_92_in_3, msg_to_check_it_14_cnu_92_in_4, msg_to_check_it_14_cnu_92_in_5, msg_to_check_it_14_cnu_93_in_0, msg_to_check_it_14_cnu_93_in_1, msg_to_check_it_14_cnu_93_in_2, msg_to_check_it_14_cnu_93_in_3, msg_to_check_it_14_cnu_93_in_4, msg_to_check_it_14_cnu_93_in_5, msg_to_check_it_14_cnu_94_in_0, msg_to_check_it_14_cnu_94_in_1, msg_to_check_it_14_cnu_94_in_2, msg_to_check_it_14_cnu_94_in_3, msg_to_check_it_14_cnu_94_in_4, msg_to_check_it_14_cnu_94_in_5, msg_to_check_it_14_cnu_95_in_0, msg_to_check_it_14_cnu_95_in_1, msg_to_check_it_14_cnu_95_in_2, msg_to_check_it_14_cnu_95_in_3, msg_to_check_it_14_cnu_95_in_4, msg_to_check_it_14_cnu_95_in_5, msg_to_check_it_14_cnu_96_in_0, msg_to_check_it_14_cnu_96_in_1, msg_to_check_it_14_cnu_96_in_2, msg_to_check_it_14_cnu_96_in_3, msg_to_check_it_14_cnu_96_in_4, msg_to_check_it_14_cnu_96_in_5, msg_to_check_it_14_cnu_97_in_0, msg_to_check_it_14_cnu_97_in_1, msg_to_check_it_14_cnu_97_in_2, msg_to_check_it_14_cnu_97_in_3, msg_to_check_it_14_cnu_97_in_4, msg_to_check_it_14_cnu_97_in_5, msg_to_check_it_14_cnu_98_in_0, msg_to_check_it_14_cnu_98_in_1, msg_to_check_it_14_cnu_98_in_2, msg_to_check_it_14_cnu_98_in_3, msg_to_check_it_14_cnu_98_in_4, msg_to_check_it_14_cnu_98_in_5, msg_to_check_it_15_cnu_0_in_0, msg_to_check_it_15_cnu_0_in_1, msg_to_check_it_15_cnu_0_in_2, msg_to_check_it_15_cnu_0_in_3, msg_to_check_it_15_cnu_0_in_4, msg_to_check_it_15_cnu_0_in_5, msg_to_check_it_15_cnu_1_in_0, msg_to_check_it_15_cnu_1_in_1, msg_to_check_it_15_cnu_1_in_2, msg_to_check_it_15_cnu_1_in_3, msg_to_check_it_15_cnu_1_in_4, msg_to_check_it_15_cnu_1_in_5, msg_to_check_it_15_cnu_2_in_0, msg_to_check_it_15_cnu_2_in_1, msg_to_check_it_15_cnu_2_in_2, msg_to_check_it_15_cnu_2_in_3, msg_to_check_it_15_cnu_2_in_4, msg_to_check_it_15_cnu_2_in_5, msg_to_check_it_15_cnu_3_in_0, msg_to_check_it_15_cnu_3_in_1, msg_to_check_it_15_cnu_3_in_2, msg_to_check_it_15_cnu_3_in_3, msg_to_check_it_15_cnu_3_in_4, msg_to_check_it_15_cnu_3_in_5, msg_to_check_it_15_cnu_4_in_0, msg_to_check_it_15_cnu_4_in_1, msg_to_check_it_15_cnu_4_in_2, msg_to_check_it_15_cnu_4_in_3, msg_to_check_it_15_cnu_4_in_4, msg_to_check_it_15_cnu_4_in_5, msg_to_check_it_15_cnu_5_in_0, msg_to_check_it_15_cnu_5_in_1, msg_to_check_it_15_cnu_5_in_2, msg_to_check_it_15_cnu_5_in_3, msg_to_check_it_15_cnu_5_in_4, msg_to_check_it_15_cnu_5_in_5, msg_to_check_it_15_cnu_6_in_0, msg_to_check_it_15_cnu_6_in_1, msg_to_check_it_15_cnu_6_in_2, msg_to_check_it_15_cnu_6_in_3, msg_to_check_it_15_cnu_6_in_4, msg_to_check_it_15_cnu_6_in_5, msg_to_check_it_15_cnu_7_in_0, msg_to_check_it_15_cnu_7_in_1, msg_to_check_it_15_cnu_7_in_2, msg_to_check_it_15_cnu_7_in_3, msg_to_check_it_15_cnu_7_in_4, msg_to_check_it_15_cnu_7_in_5, msg_to_check_it_15_cnu_8_in_0, msg_to_check_it_15_cnu_8_in_1, msg_to_check_it_15_cnu_8_in_2, msg_to_check_it_15_cnu_8_in_3, msg_to_check_it_15_cnu_8_in_4, msg_to_check_it_15_cnu_8_in_5, msg_to_check_it_15_cnu_9_in_0, msg_to_check_it_15_cnu_9_in_1, msg_to_check_it_15_cnu_9_in_2, msg_to_check_it_15_cnu_9_in_3, msg_to_check_it_15_cnu_9_in_4, msg_to_check_it_15_cnu_9_in_5, msg_to_check_it_15_cnu_10_in_0, msg_to_check_it_15_cnu_10_in_1, msg_to_check_it_15_cnu_10_in_2, msg_to_check_it_15_cnu_10_in_3, msg_to_check_it_15_cnu_10_in_4, msg_to_check_it_15_cnu_10_in_5, msg_to_check_it_15_cnu_11_in_0, msg_to_check_it_15_cnu_11_in_1, msg_to_check_it_15_cnu_11_in_2, msg_to_check_it_15_cnu_11_in_3, msg_to_check_it_15_cnu_11_in_4, msg_to_check_it_15_cnu_11_in_5, msg_to_check_it_15_cnu_12_in_0, msg_to_check_it_15_cnu_12_in_1, msg_to_check_it_15_cnu_12_in_2, msg_to_check_it_15_cnu_12_in_3, msg_to_check_it_15_cnu_12_in_4, msg_to_check_it_15_cnu_12_in_5, msg_to_check_it_15_cnu_13_in_0, msg_to_check_it_15_cnu_13_in_1, msg_to_check_it_15_cnu_13_in_2, msg_to_check_it_15_cnu_13_in_3, msg_to_check_it_15_cnu_13_in_4, msg_to_check_it_15_cnu_13_in_5, msg_to_check_it_15_cnu_14_in_0, msg_to_check_it_15_cnu_14_in_1, msg_to_check_it_15_cnu_14_in_2, msg_to_check_it_15_cnu_14_in_3, msg_to_check_it_15_cnu_14_in_4, msg_to_check_it_15_cnu_14_in_5, msg_to_check_it_15_cnu_15_in_0, msg_to_check_it_15_cnu_15_in_1, msg_to_check_it_15_cnu_15_in_2, msg_to_check_it_15_cnu_15_in_3, msg_to_check_it_15_cnu_15_in_4, msg_to_check_it_15_cnu_15_in_5, msg_to_check_it_15_cnu_16_in_0, msg_to_check_it_15_cnu_16_in_1, msg_to_check_it_15_cnu_16_in_2, msg_to_check_it_15_cnu_16_in_3, msg_to_check_it_15_cnu_16_in_4, msg_to_check_it_15_cnu_16_in_5, msg_to_check_it_15_cnu_17_in_0, msg_to_check_it_15_cnu_17_in_1, msg_to_check_it_15_cnu_17_in_2, msg_to_check_it_15_cnu_17_in_3, msg_to_check_it_15_cnu_17_in_4, msg_to_check_it_15_cnu_17_in_5, msg_to_check_it_15_cnu_18_in_0, msg_to_check_it_15_cnu_18_in_1, msg_to_check_it_15_cnu_18_in_2, msg_to_check_it_15_cnu_18_in_3, msg_to_check_it_15_cnu_18_in_4, msg_to_check_it_15_cnu_18_in_5, msg_to_check_it_15_cnu_19_in_0, msg_to_check_it_15_cnu_19_in_1, msg_to_check_it_15_cnu_19_in_2, msg_to_check_it_15_cnu_19_in_3, msg_to_check_it_15_cnu_19_in_4, msg_to_check_it_15_cnu_19_in_5, msg_to_check_it_15_cnu_20_in_0, msg_to_check_it_15_cnu_20_in_1, msg_to_check_it_15_cnu_20_in_2, msg_to_check_it_15_cnu_20_in_3, msg_to_check_it_15_cnu_20_in_4, msg_to_check_it_15_cnu_20_in_5, msg_to_check_it_15_cnu_21_in_0, msg_to_check_it_15_cnu_21_in_1, msg_to_check_it_15_cnu_21_in_2, msg_to_check_it_15_cnu_21_in_3, msg_to_check_it_15_cnu_21_in_4, msg_to_check_it_15_cnu_21_in_5, msg_to_check_it_15_cnu_22_in_0, msg_to_check_it_15_cnu_22_in_1, msg_to_check_it_15_cnu_22_in_2, msg_to_check_it_15_cnu_22_in_3, msg_to_check_it_15_cnu_22_in_4, msg_to_check_it_15_cnu_22_in_5, msg_to_check_it_15_cnu_23_in_0, msg_to_check_it_15_cnu_23_in_1, msg_to_check_it_15_cnu_23_in_2, msg_to_check_it_15_cnu_23_in_3, msg_to_check_it_15_cnu_23_in_4, msg_to_check_it_15_cnu_23_in_5, msg_to_check_it_15_cnu_24_in_0, msg_to_check_it_15_cnu_24_in_1, msg_to_check_it_15_cnu_24_in_2, msg_to_check_it_15_cnu_24_in_3, msg_to_check_it_15_cnu_24_in_4, msg_to_check_it_15_cnu_24_in_5, msg_to_check_it_15_cnu_25_in_0, msg_to_check_it_15_cnu_25_in_1, msg_to_check_it_15_cnu_25_in_2, msg_to_check_it_15_cnu_25_in_3, msg_to_check_it_15_cnu_25_in_4, msg_to_check_it_15_cnu_25_in_5, msg_to_check_it_15_cnu_26_in_0, msg_to_check_it_15_cnu_26_in_1, msg_to_check_it_15_cnu_26_in_2, msg_to_check_it_15_cnu_26_in_3, msg_to_check_it_15_cnu_26_in_4, msg_to_check_it_15_cnu_26_in_5, msg_to_check_it_15_cnu_27_in_0, msg_to_check_it_15_cnu_27_in_1, msg_to_check_it_15_cnu_27_in_2, msg_to_check_it_15_cnu_27_in_3, msg_to_check_it_15_cnu_27_in_4, msg_to_check_it_15_cnu_27_in_5, msg_to_check_it_15_cnu_28_in_0, msg_to_check_it_15_cnu_28_in_1, msg_to_check_it_15_cnu_28_in_2, msg_to_check_it_15_cnu_28_in_3, msg_to_check_it_15_cnu_28_in_4, msg_to_check_it_15_cnu_28_in_5, msg_to_check_it_15_cnu_29_in_0, msg_to_check_it_15_cnu_29_in_1, msg_to_check_it_15_cnu_29_in_2, msg_to_check_it_15_cnu_29_in_3, msg_to_check_it_15_cnu_29_in_4, msg_to_check_it_15_cnu_29_in_5, msg_to_check_it_15_cnu_30_in_0, msg_to_check_it_15_cnu_30_in_1, msg_to_check_it_15_cnu_30_in_2, msg_to_check_it_15_cnu_30_in_3, msg_to_check_it_15_cnu_30_in_4, msg_to_check_it_15_cnu_30_in_5, msg_to_check_it_15_cnu_31_in_0, msg_to_check_it_15_cnu_31_in_1, msg_to_check_it_15_cnu_31_in_2, msg_to_check_it_15_cnu_31_in_3, msg_to_check_it_15_cnu_31_in_4, msg_to_check_it_15_cnu_31_in_5, msg_to_check_it_15_cnu_32_in_0, msg_to_check_it_15_cnu_32_in_1, msg_to_check_it_15_cnu_32_in_2, msg_to_check_it_15_cnu_32_in_3, msg_to_check_it_15_cnu_32_in_4, msg_to_check_it_15_cnu_32_in_5, msg_to_check_it_15_cnu_33_in_0, msg_to_check_it_15_cnu_33_in_1, msg_to_check_it_15_cnu_33_in_2, msg_to_check_it_15_cnu_33_in_3, msg_to_check_it_15_cnu_33_in_4, msg_to_check_it_15_cnu_33_in_5, msg_to_check_it_15_cnu_34_in_0, msg_to_check_it_15_cnu_34_in_1, msg_to_check_it_15_cnu_34_in_2, msg_to_check_it_15_cnu_34_in_3, msg_to_check_it_15_cnu_34_in_4, msg_to_check_it_15_cnu_34_in_5, msg_to_check_it_15_cnu_35_in_0, msg_to_check_it_15_cnu_35_in_1, msg_to_check_it_15_cnu_35_in_2, msg_to_check_it_15_cnu_35_in_3, msg_to_check_it_15_cnu_35_in_4, msg_to_check_it_15_cnu_35_in_5, msg_to_check_it_15_cnu_36_in_0, msg_to_check_it_15_cnu_36_in_1, msg_to_check_it_15_cnu_36_in_2, msg_to_check_it_15_cnu_36_in_3, msg_to_check_it_15_cnu_36_in_4, msg_to_check_it_15_cnu_36_in_5, msg_to_check_it_15_cnu_37_in_0, msg_to_check_it_15_cnu_37_in_1, msg_to_check_it_15_cnu_37_in_2, msg_to_check_it_15_cnu_37_in_3, msg_to_check_it_15_cnu_37_in_4, msg_to_check_it_15_cnu_37_in_5, msg_to_check_it_15_cnu_38_in_0, msg_to_check_it_15_cnu_38_in_1, msg_to_check_it_15_cnu_38_in_2, msg_to_check_it_15_cnu_38_in_3, msg_to_check_it_15_cnu_38_in_4, msg_to_check_it_15_cnu_38_in_5, msg_to_check_it_15_cnu_39_in_0, msg_to_check_it_15_cnu_39_in_1, msg_to_check_it_15_cnu_39_in_2, msg_to_check_it_15_cnu_39_in_3, msg_to_check_it_15_cnu_39_in_4, msg_to_check_it_15_cnu_39_in_5, msg_to_check_it_15_cnu_40_in_0, msg_to_check_it_15_cnu_40_in_1, msg_to_check_it_15_cnu_40_in_2, msg_to_check_it_15_cnu_40_in_3, msg_to_check_it_15_cnu_40_in_4, msg_to_check_it_15_cnu_40_in_5, msg_to_check_it_15_cnu_41_in_0, msg_to_check_it_15_cnu_41_in_1, msg_to_check_it_15_cnu_41_in_2, msg_to_check_it_15_cnu_41_in_3, msg_to_check_it_15_cnu_41_in_4, msg_to_check_it_15_cnu_41_in_5, msg_to_check_it_15_cnu_42_in_0, msg_to_check_it_15_cnu_42_in_1, msg_to_check_it_15_cnu_42_in_2, msg_to_check_it_15_cnu_42_in_3, msg_to_check_it_15_cnu_42_in_4, msg_to_check_it_15_cnu_42_in_5, msg_to_check_it_15_cnu_43_in_0, msg_to_check_it_15_cnu_43_in_1, msg_to_check_it_15_cnu_43_in_2, msg_to_check_it_15_cnu_43_in_3, msg_to_check_it_15_cnu_43_in_4, msg_to_check_it_15_cnu_43_in_5, msg_to_check_it_15_cnu_44_in_0, msg_to_check_it_15_cnu_44_in_1, msg_to_check_it_15_cnu_44_in_2, msg_to_check_it_15_cnu_44_in_3, msg_to_check_it_15_cnu_44_in_4, msg_to_check_it_15_cnu_44_in_5, msg_to_check_it_15_cnu_45_in_0, msg_to_check_it_15_cnu_45_in_1, msg_to_check_it_15_cnu_45_in_2, msg_to_check_it_15_cnu_45_in_3, msg_to_check_it_15_cnu_45_in_4, msg_to_check_it_15_cnu_45_in_5, msg_to_check_it_15_cnu_46_in_0, msg_to_check_it_15_cnu_46_in_1, msg_to_check_it_15_cnu_46_in_2, msg_to_check_it_15_cnu_46_in_3, msg_to_check_it_15_cnu_46_in_4, msg_to_check_it_15_cnu_46_in_5, msg_to_check_it_15_cnu_47_in_0, msg_to_check_it_15_cnu_47_in_1, msg_to_check_it_15_cnu_47_in_2, msg_to_check_it_15_cnu_47_in_3, msg_to_check_it_15_cnu_47_in_4, msg_to_check_it_15_cnu_47_in_5, msg_to_check_it_15_cnu_48_in_0, msg_to_check_it_15_cnu_48_in_1, msg_to_check_it_15_cnu_48_in_2, msg_to_check_it_15_cnu_48_in_3, msg_to_check_it_15_cnu_48_in_4, msg_to_check_it_15_cnu_48_in_5, msg_to_check_it_15_cnu_49_in_0, msg_to_check_it_15_cnu_49_in_1, msg_to_check_it_15_cnu_49_in_2, msg_to_check_it_15_cnu_49_in_3, msg_to_check_it_15_cnu_49_in_4, msg_to_check_it_15_cnu_49_in_5, msg_to_check_it_15_cnu_50_in_0, msg_to_check_it_15_cnu_50_in_1, msg_to_check_it_15_cnu_50_in_2, msg_to_check_it_15_cnu_50_in_3, msg_to_check_it_15_cnu_50_in_4, msg_to_check_it_15_cnu_50_in_5, msg_to_check_it_15_cnu_51_in_0, msg_to_check_it_15_cnu_51_in_1, msg_to_check_it_15_cnu_51_in_2, msg_to_check_it_15_cnu_51_in_3, msg_to_check_it_15_cnu_51_in_4, msg_to_check_it_15_cnu_51_in_5, msg_to_check_it_15_cnu_52_in_0, msg_to_check_it_15_cnu_52_in_1, msg_to_check_it_15_cnu_52_in_2, msg_to_check_it_15_cnu_52_in_3, msg_to_check_it_15_cnu_52_in_4, msg_to_check_it_15_cnu_52_in_5, msg_to_check_it_15_cnu_53_in_0, msg_to_check_it_15_cnu_53_in_1, msg_to_check_it_15_cnu_53_in_2, msg_to_check_it_15_cnu_53_in_3, msg_to_check_it_15_cnu_53_in_4, msg_to_check_it_15_cnu_53_in_5, msg_to_check_it_15_cnu_54_in_0, msg_to_check_it_15_cnu_54_in_1, msg_to_check_it_15_cnu_54_in_2, msg_to_check_it_15_cnu_54_in_3, msg_to_check_it_15_cnu_54_in_4, msg_to_check_it_15_cnu_54_in_5, msg_to_check_it_15_cnu_55_in_0, msg_to_check_it_15_cnu_55_in_1, msg_to_check_it_15_cnu_55_in_2, msg_to_check_it_15_cnu_55_in_3, msg_to_check_it_15_cnu_55_in_4, msg_to_check_it_15_cnu_55_in_5, msg_to_check_it_15_cnu_56_in_0, msg_to_check_it_15_cnu_56_in_1, msg_to_check_it_15_cnu_56_in_2, msg_to_check_it_15_cnu_56_in_3, msg_to_check_it_15_cnu_56_in_4, msg_to_check_it_15_cnu_56_in_5, msg_to_check_it_15_cnu_57_in_0, msg_to_check_it_15_cnu_57_in_1, msg_to_check_it_15_cnu_57_in_2, msg_to_check_it_15_cnu_57_in_3, msg_to_check_it_15_cnu_57_in_4, msg_to_check_it_15_cnu_57_in_5, msg_to_check_it_15_cnu_58_in_0, msg_to_check_it_15_cnu_58_in_1, msg_to_check_it_15_cnu_58_in_2, msg_to_check_it_15_cnu_58_in_3, msg_to_check_it_15_cnu_58_in_4, msg_to_check_it_15_cnu_58_in_5, msg_to_check_it_15_cnu_59_in_0, msg_to_check_it_15_cnu_59_in_1, msg_to_check_it_15_cnu_59_in_2, msg_to_check_it_15_cnu_59_in_3, msg_to_check_it_15_cnu_59_in_4, msg_to_check_it_15_cnu_59_in_5, msg_to_check_it_15_cnu_60_in_0, msg_to_check_it_15_cnu_60_in_1, msg_to_check_it_15_cnu_60_in_2, msg_to_check_it_15_cnu_60_in_3, msg_to_check_it_15_cnu_60_in_4, msg_to_check_it_15_cnu_60_in_5, msg_to_check_it_15_cnu_61_in_0, msg_to_check_it_15_cnu_61_in_1, msg_to_check_it_15_cnu_61_in_2, msg_to_check_it_15_cnu_61_in_3, msg_to_check_it_15_cnu_61_in_4, msg_to_check_it_15_cnu_61_in_5, msg_to_check_it_15_cnu_62_in_0, msg_to_check_it_15_cnu_62_in_1, msg_to_check_it_15_cnu_62_in_2, msg_to_check_it_15_cnu_62_in_3, msg_to_check_it_15_cnu_62_in_4, msg_to_check_it_15_cnu_62_in_5, msg_to_check_it_15_cnu_63_in_0, msg_to_check_it_15_cnu_63_in_1, msg_to_check_it_15_cnu_63_in_2, msg_to_check_it_15_cnu_63_in_3, msg_to_check_it_15_cnu_63_in_4, msg_to_check_it_15_cnu_63_in_5, msg_to_check_it_15_cnu_64_in_0, msg_to_check_it_15_cnu_64_in_1, msg_to_check_it_15_cnu_64_in_2, msg_to_check_it_15_cnu_64_in_3, msg_to_check_it_15_cnu_64_in_4, msg_to_check_it_15_cnu_64_in_5, msg_to_check_it_15_cnu_65_in_0, msg_to_check_it_15_cnu_65_in_1, msg_to_check_it_15_cnu_65_in_2, msg_to_check_it_15_cnu_65_in_3, msg_to_check_it_15_cnu_65_in_4, msg_to_check_it_15_cnu_65_in_5, msg_to_check_it_15_cnu_66_in_0, msg_to_check_it_15_cnu_66_in_1, msg_to_check_it_15_cnu_66_in_2, msg_to_check_it_15_cnu_66_in_3, msg_to_check_it_15_cnu_66_in_4, msg_to_check_it_15_cnu_66_in_5, msg_to_check_it_15_cnu_67_in_0, msg_to_check_it_15_cnu_67_in_1, msg_to_check_it_15_cnu_67_in_2, msg_to_check_it_15_cnu_67_in_3, msg_to_check_it_15_cnu_67_in_4, msg_to_check_it_15_cnu_67_in_5, msg_to_check_it_15_cnu_68_in_0, msg_to_check_it_15_cnu_68_in_1, msg_to_check_it_15_cnu_68_in_2, msg_to_check_it_15_cnu_68_in_3, msg_to_check_it_15_cnu_68_in_4, msg_to_check_it_15_cnu_68_in_5, msg_to_check_it_15_cnu_69_in_0, msg_to_check_it_15_cnu_69_in_1, msg_to_check_it_15_cnu_69_in_2, msg_to_check_it_15_cnu_69_in_3, msg_to_check_it_15_cnu_69_in_4, msg_to_check_it_15_cnu_69_in_5, msg_to_check_it_15_cnu_70_in_0, msg_to_check_it_15_cnu_70_in_1, msg_to_check_it_15_cnu_70_in_2, msg_to_check_it_15_cnu_70_in_3, msg_to_check_it_15_cnu_70_in_4, msg_to_check_it_15_cnu_70_in_5, msg_to_check_it_15_cnu_71_in_0, msg_to_check_it_15_cnu_71_in_1, msg_to_check_it_15_cnu_71_in_2, msg_to_check_it_15_cnu_71_in_3, msg_to_check_it_15_cnu_71_in_4, msg_to_check_it_15_cnu_71_in_5, msg_to_check_it_15_cnu_72_in_0, msg_to_check_it_15_cnu_72_in_1, msg_to_check_it_15_cnu_72_in_2, msg_to_check_it_15_cnu_72_in_3, msg_to_check_it_15_cnu_72_in_4, msg_to_check_it_15_cnu_72_in_5, msg_to_check_it_15_cnu_73_in_0, msg_to_check_it_15_cnu_73_in_1, msg_to_check_it_15_cnu_73_in_2, msg_to_check_it_15_cnu_73_in_3, msg_to_check_it_15_cnu_73_in_4, msg_to_check_it_15_cnu_73_in_5, msg_to_check_it_15_cnu_74_in_0, msg_to_check_it_15_cnu_74_in_1, msg_to_check_it_15_cnu_74_in_2, msg_to_check_it_15_cnu_74_in_3, msg_to_check_it_15_cnu_74_in_4, msg_to_check_it_15_cnu_74_in_5, msg_to_check_it_15_cnu_75_in_0, msg_to_check_it_15_cnu_75_in_1, msg_to_check_it_15_cnu_75_in_2, msg_to_check_it_15_cnu_75_in_3, msg_to_check_it_15_cnu_75_in_4, msg_to_check_it_15_cnu_75_in_5, msg_to_check_it_15_cnu_76_in_0, msg_to_check_it_15_cnu_76_in_1, msg_to_check_it_15_cnu_76_in_2, msg_to_check_it_15_cnu_76_in_3, msg_to_check_it_15_cnu_76_in_4, msg_to_check_it_15_cnu_76_in_5, msg_to_check_it_15_cnu_77_in_0, msg_to_check_it_15_cnu_77_in_1, msg_to_check_it_15_cnu_77_in_2, msg_to_check_it_15_cnu_77_in_3, msg_to_check_it_15_cnu_77_in_4, msg_to_check_it_15_cnu_77_in_5, msg_to_check_it_15_cnu_78_in_0, msg_to_check_it_15_cnu_78_in_1, msg_to_check_it_15_cnu_78_in_2, msg_to_check_it_15_cnu_78_in_3, msg_to_check_it_15_cnu_78_in_4, msg_to_check_it_15_cnu_78_in_5, msg_to_check_it_15_cnu_79_in_0, msg_to_check_it_15_cnu_79_in_1, msg_to_check_it_15_cnu_79_in_2, msg_to_check_it_15_cnu_79_in_3, msg_to_check_it_15_cnu_79_in_4, msg_to_check_it_15_cnu_79_in_5, msg_to_check_it_15_cnu_80_in_0, msg_to_check_it_15_cnu_80_in_1, msg_to_check_it_15_cnu_80_in_2, msg_to_check_it_15_cnu_80_in_3, msg_to_check_it_15_cnu_80_in_4, msg_to_check_it_15_cnu_80_in_5, msg_to_check_it_15_cnu_81_in_0, msg_to_check_it_15_cnu_81_in_1, msg_to_check_it_15_cnu_81_in_2, msg_to_check_it_15_cnu_81_in_3, msg_to_check_it_15_cnu_81_in_4, msg_to_check_it_15_cnu_81_in_5, msg_to_check_it_15_cnu_82_in_0, msg_to_check_it_15_cnu_82_in_1, msg_to_check_it_15_cnu_82_in_2, msg_to_check_it_15_cnu_82_in_3, msg_to_check_it_15_cnu_82_in_4, msg_to_check_it_15_cnu_82_in_5, msg_to_check_it_15_cnu_83_in_0, msg_to_check_it_15_cnu_83_in_1, msg_to_check_it_15_cnu_83_in_2, msg_to_check_it_15_cnu_83_in_3, msg_to_check_it_15_cnu_83_in_4, msg_to_check_it_15_cnu_83_in_5, msg_to_check_it_15_cnu_84_in_0, msg_to_check_it_15_cnu_84_in_1, msg_to_check_it_15_cnu_84_in_2, msg_to_check_it_15_cnu_84_in_3, msg_to_check_it_15_cnu_84_in_4, msg_to_check_it_15_cnu_84_in_5, msg_to_check_it_15_cnu_85_in_0, msg_to_check_it_15_cnu_85_in_1, msg_to_check_it_15_cnu_85_in_2, msg_to_check_it_15_cnu_85_in_3, msg_to_check_it_15_cnu_85_in_4, msg_to_check_it_15_cnu_85_in_5, msg_to_check_it_15_cnu_86_in_0, msg_to_check_it_15_cnu_86_in_1, msg_to_check_it_15_cnu_86_in_2, msg_to_check_it_15_cnu_86_in_3, msg_to_check_it_15_cnu_86_in_4, msg_to_check_it_15_cnu_86_in_5, msg_to_check_it_15_cnu_87_in_0, msg_to_check_it_15_cnu_87_in_1, msg_to_check_it_15_cnu_87_in_2, msg_to_check_it_15_cnu_87_in_3, msg_to_check_it_15_cnu_87_in_4, msg_to_check_it_15_cnu_87_in_5, msg_to_check_it_15_cnu_88_in_0, msg_to_check_it_15_cnu_88_in_1, msg_to_check_it_15_cnu_88_in_2, msg_to_check_it_15_cnu_88_in_3, msg_to_check_it_15_cnu_88_in_4, msg_to_check_it_15_cnu_88_in_5, msg_to_check_it_15_cnu_89_in_0, msg_to_check_it_15_cnu_89_in_1, msg_to_check_it_15_cnu_89_in_2, msg_to_check_it_15_cnu_89_in_3, msg_to_check_it_15_cnu_89_in_4, msg_to_check_it_15_cnu_89_in_5, msg_to_check_it_15_cnu_90_in_0, msg_to_check_it_15_cnu_90_in_1, msg_to_check_it_15_cnu_90_in_2, msg_to_check_it_15_cnu_90_in_3, msg_to_check_it_15_cnu_90_in_4, msg_to_check_it_15_cnu_90_in_5, msg_to_check_it_15_cnu_91_in_0, msg_to_check_it_15_cnu_91_in_1, msg_to_check_it_15_cnu_91_in_2, msg_to_check_it_15_cnu_91_in_3, msg_to_check_it_15_cnu_91_in_4, msg_to_check_it_15_cnu_91_in_5, msg_to_check_it_15_cnu_92_in_0, msg_to_check_it_15_cnu_92_in_1, msg_to_check_it_15_cnu_92_in_2, msg_to_check_it_15_cnu_92_in_3, msg_to_check_it_15_cnu_92_in_4, msg_to_check_it_15_cnu_92_in_5, msg_to_check_it_15_cnu_93_in_0, msg_to_check_it_15_cnu_93_in_1, msg_to_check_it_15_cnu_93_in_2, msg_to_check_it_15_cnu_93_in_3, msg_to_check_it_15_cnu_93_in_4, msg_to_check_it_15_cnu_93_in_5, msg_to_check_it_15_cnu_94_in_0, msg_to_check_it_15_cnu_94_in_1, msg_to_check_it_15_cnu_94_in_2, msg_to_check_it_15_cnu_94_in_3, msg_to_check_it_15_cnu_94_in_4, msg_to_check_it_15_cnu_94_in_5, msg_to_check_it_15_cnu_95_in_0, msg_to_check_it_15_cnu_95_in_1, msg_to_check_it_15_cnu_95_in_2, msg_to_check_it_15_cnu_95_in_3, msg_to_check_it_15_cnu_95_in_4, msg_to_check_it_15_cnu_95_in_5, msg_to_check_it_15_cnu_96_in_0, msg_to_check_it_15_cnu_96_in_1, msg_to_check_it_15_cnu_96_in_2, msg_to_check_it_15_cnu_96_in_3, msg_to_check_it_15_cnu_96_in_4, msg_to_check_it_15_cnu_96_in_5, msg_to_check_it_15_cnu_97_in_0, msg_to_check_it_15_cnu_97_in_1, msg_to_check_it_15_cnu_97_in_2, msg_to_check_it_15_cnu_97_in_3, msg_to_check_it_15_cnu_97_in_4, msg_to_check_it_15_cnu_97_in_5, msg_to_check_it_15_cnu_98_in_0, msg_to_check_it_15_cnu_98_in_1, msg_to_check_it_15_cnu_98_in_2, msg_to_check_it_15_cnu_98_in_3, msg_to_check_it_15_cnu_98_in_4, msg_to_check_it_15_cnu_98_in_5, msg_to_check_it_16_cnu_0_in_0, msg_to_check_it_16_cnu_0_in_1, msg_to_check_it_16_cnu_0_in_2, msg_to_check_it_16_cnu_0_in_3, msg_to_check_it_16_cnu_0_in_4, msg_to_check_it_16_cnu_0_in_5, msg_to_check_it_16_cnu_1_in_0, msg_to_check_it_16_cnu_1_in_1, msg_to_check_it_16_cnu_1_in_2, msg_to_check_it_16_cnu_1_in_3, msg_to_check_it_16_cnu_1_in_4, msg_to_check_it_16_cnu_1_in_5, msg_to_check_it_16_cnu_2_in_0, msg_to_check_it_16_cnu_2_in_1, msg_to_check_it_16_cnu_2_in_2, msg_to_check_it_16_cnu_2_in_3, msg_to_check_it_16_cnu_2_in_4, msg_to_check_it_16_cnu_2_in_5, msg_to_check_it_16_cnu_3_in_0, msg_to_check_it_16_cnu_3_in_1, msg_to_check_it_16_cnu_3_in_2, msg_to_check_it_16_cnu_3_in_3, msg_to_check_it_16_cnu_3_in_4, msg_to_check_it_16_cnu_3_in_5, msg_to_check_it_16_cnu_4_in_0, msg_to_check_it_16_cnu_4_in_1, msg_to_check_it_16_cnu_4_in_2, msg_to_check_it_16_cnu_4_in_3, msg_to_check_it_16_cnu_4_in_4, msg_to_check_it_16_cnu_4_in_5, msg_to_check_it_16_cnu_5_in_0, msg_to_check_it_16_cnu_5_in_1, msg_to_check_it_16_cnu_5_in_2, msg_to_check_it_16_cnu_5_in_3, msg_to_check_it_16_cnu_5_in_4, msg_to_check_it_16_cnu_5_in_5, msg_to_check_it_16_cnu_6_in_0, msg_to_check_it_16_cnu_6_in_1, msg_to_check_it_16_cnu_6_in_2, msg_to_check_it_16_cnu_6_in_3, msg_to_check_it_16_cnu_6_in_4, msg_to_check_it_16_cnu_6_in_5, msg_to_check_it_16_cnu_7_in_0, msg_to_check_it_16_cnu_7_in_1, msg_to_check_it_16_cnu_7_in_2, msg_to_check_it_16_cnu_7_in_3, msg_to_check_it_16_cnu_7_in_4, msg_to_check_it_16_cnu_7_in_5, msg_to_check_it_16_cnu_8_in_0, msg_to_check_it_16_cnu_8_in_1, msg_to_check_it_16_cnu_8_in_2, msg_to_check_it_16_cnu_8_in_3, msg_to_check_it_16_cnu_8_in_4, msg_to_check_it_16_cnu_8_in_5, msg_to_check_it_16_cnu_9_in_0, msg_to_check_it_16_cnu_9_in_1, msg_to_check_it_16_cnu_9_in_2, msg_to_check_it_16_cnu_9_in_3, msg_to_check_it_16_cnu_9_in_4, msg_to_check_it_16_cnu_9_in_5, msg_to_check_it_16_cnu_10_in_0, msg_to_check_it_16_cnu_10_in_1, msg_to_check_it_16_cnu_10_in_2, msg_to_check_it_16_cnu_10_in_3, msg_to_check_it_16_cnu_10_in_4, msg_to_check_it_16_cnu_10_in_5, msg_to_check_it_16_cnu_11_in_0, msg_to_check_it_16_cnu_11_in_1, msg_to_check_it_16_cnu_11_in_2, msg_to_check_it_16_cnu_11_in_3, msg_to_check_it_16_cnu_11_in_4, msg_to_check_it_16_cnu_11_in_5, msg_to_check_it_16_cnu_12_in_0, msg_to_check_it_16_cnu_12_in_1, msg_to_check_it_16_cnu_12_in_2, msg_to_check_it_16_cnu_12_in_3, msg_to_check_it_16_cnu_12_in_4, msg_to_check_it_16_cnu_12_in_5, msg_to_check_it_16_cnu_13_in_0, msg_to_check_it_16_cnu_13_in_1, msg_to_check_it_16_cnu_13_in_2, msg_to_check_it_16_cnu_13_in_3, msg_to_check_it_16_cnu_13_in_4, msg_to_check_it_16_cnu_13_in_5, msg_to_check_it_16_cnu_14_in_0, msg_to_check_it_16_cnu_14_in_1, msg_to_check_it_16_cnu_14_in_2, msg_to_check_it_16_cnu_14_in_3, msg_to_check_it_16_cnu_14_in_4, msg_to_check_it_16_cnu_14_in_5, msg_to_check_it_16_cnu_15_in_0, msg_to_check_it_16_cnu_15_in_1, msg_to_check_it_16_cnu_15_in_2, msg_to_check_it_16_cnu_15_in_3, msg_to_check_it_16_cnu_15_in_4, msg_to_check_it_16_cnu_15_in_5, msg_to_check_it_16_cnu_16_in_0, msg_to_check_it_16_cnu_16_in_1, msg_to_check_it_16_cnu_16_in_2, msg_to_check_it_16_cnu_16_in_3, msg_to_check_it_16_cnu_16_in_4, msg_to_check_it_16_cnu_16_in_5, msg_to_check_it_16_cnu_17_in_0, msg_to_check_it_16_cnu_17_in_1, msg_to_check_it_16_cnu_17_in_2, msg_to_check_it_16_cnu_17_in_3, msg_to_check_it_16_cnu_17_in_4, msg_to_check_it_16_cnu_17_in_5, msg_to_check_it_16_cnu_18_in_0, msg_to_check_it_16_cnu_18_in_1, msg_to_check_it_16_cnu_18_in_2, msg_to_check_it_16_cnu_18_in_3, msg_to_check_it_16_cnu_18_in_4, msg_to_check_it_16_cnu_18_in_5, msg_to_check_it_16_cnu_19_in_0, msg_to_check_it_16_cnu_19_in_1, msg_to_check_it_16_cnu_19_in_2, msg_to_check_it_16_cnu_19_in_3, msg_to_check_it_16_cnu_19_in_4, msg_to_check_it_16_cnu_19_in_5, msg_to_check_it_16_cnu_20_in_0, msg_to_check_it_16_cnu_20_in_1, msg_to_check_it_16_cnu_20_in_2, msg_to_check_it_16_cnu_20_in_3, msg_to_check_it_16_cnu_20_in_4, msg_to_check_it_16_cnu_20_in_5, msg_to_check_it_16_cnu_21_in_0, msg_to_check_it_16_cnu_21_in_1, msg_to_check_it_16_cnu_21_in_2, msg_to_check_it_16_cnu_21_in_3, msg_to_check_it_16_cnu_21_in_4, msg_to_check_it_16_cnu_21_in_5, msg_to_check_it_16_cnu_22_in_0, msg_to_check_it_16_cnu_22_in_1, msg_to_check_it_16_cnu_22_in_2, msg_to_check_it_16_cnu_22_in_3, msg_to_check_it_16_cnu_22_in_4, msg_to_check_it_16_cnu_22_in_5, msg_to_check_it_16_cnu_23_in_0, msg_to_check_it_16_cnu_23_in_1, msg_to_check_it_16_cnu_23_in_2, msg_to_check_it_16_cnu_23_in_3, msg_to_check_it_16_cnu_23_in_4, msg_to_check_it_16_cnu_23_in_5, msg_to_check_it_16_cnu_24_in_0, msg_to_check_it_16_cnu_24_in_1, msg_to_check_it_16_cnu_24_in_2, msg_to_check_it_16_cnu_24_in_3, msg_to_check_it_16_cnu_24_in_4, msg_to_check_it_16_cnu_24_in_5, msg_to_check_it_16_cnu_25_in_0, msg_to_check_it_16_cnu_25_in_1, msg_to_check_it_16_cnu_25_in_2, msg_to_check_it_16_cnu_25_in_3, msg_to_check_it_16_cnu_25_in_4, msg_to_check_it_16_cnu_25_in_5, msg_to_check_it_16_cnu_26_in_0, msg_to_check_it_16_cnu_26_in_1, msg_to_check_it_16_cnu_26_in_2, msg_to_check_it_16_cnu_26_in_3, msg_to_check_it_16_cnu_26_in_4, msg_to_check_it_16_cnu_26_in_5, msg_to_check_it_16_cnu_27_in_0, msg_to_check_it_16_cnu_27_in_1, msg_to_check_it_16_cnu_27_in_2, msg_to_check_it_16_cnu_27_in_3, msg_to_check_it_16_cnu_27_in_4, msg_to_check_it_16_cnu_27_in_5, msg_to_check_it_16_cnu_28_in_0, msg_to_check_it_16_cnu_28_in_1, msg_to_check_it_16_cnu_28_in_2, msg_to_check_it_16_cnu_28_in_3, msg_to_check_it_16_cnu_28_in_4, msg_to_check_it_16_cnu_28_in_5, msg_to_check_it_16_cnu_29_in_0, msg_to_check_it_16_cnu_29_in_1, msg_to_check_it_16_cnu_29_in_2, msg_to_check_it_16_cnu_29_in_3, msg_to_check_it_16_cnu_29_in_4, msg_to_check_it_16_cnu_29_in_5, msg_to_check_it_16_cnu_30_in_0, msg_to_check_it_16_cnu_30_in_1, msg_to_check_it_16_cnu_30_in_2, msg_to_check_it_16_cnu_30_in_3, msg_to_check_it_16_cnu_30_in_4, msg_to_check_it_16_cnu_30_in_5, msg_to_check_it_16_cnu_31_in_0, msg_to_check_it_16_cnu_31_in_1, msg_to_check_it_16_cnu_31_in_2, msg_to_check_it_16_cnu_31_in_3, msg_to_check_it_16_cnu_31_in_4, msg_to_check_it_16_cnu_31_in_5, msg_to_check_it_16_cnu_32_in_0, msg_to_check_it_16_cnu_32_in_1, msg_to_check_it_16_cnu_32_in_2, msg_to_check_it_16_cnu_32_in_3, msg_to_check_it_16_cnu_32_in_4, msg_to_check_it_16_cnu_32_in_5, msg_to_check_it_16_cnu_33_in_0, msg_to_check_it_16_cnu_33_in_1, msg_to_check_it_16_cnu_33_in_2, msg_to_check_it_16_cnu_33_in_3, msg_to_check_it_16_cnu_33_in_4, msg_to_check_it_16_cnu_33_in_5, msg_to_check_it_16_cnu_34_in_0, msg_to_check_it_16_cnu_34_in_1, msg_to_check_it_16_cnu_34_in_2, msg_to_check_it_16_cnu_34_in_3, msg_to_check_it_16_cnu_34_in_4, msg_to_check_it_16_cnu_34_in_5, msg_to_check_it_16_cnu_35_in_0, msg_to_check_it_16_cnu_35_in_1, msg_to_check_it_16_cnu_35_in_2, msg_to_check_it_16_cnu_35_in_3, msg_to_check_it_16_cnu_35_in_4, msg_to_check_it_16_cnu_35_in_5, msg_to_check_it_16_cnu_36_in_0, msg_to_check_it_16_cnu_36_in_1, msg_to_check_it_16_cnu_36_in_2, msg_to_check_it_16_cnu_36_in_3, msg_to_check_it_16_cnu_36_in_4, msg_to_check_it_16_cnu_36_in_5, msg_to_check_it_16_cnu_37_in_0, msg_to_check_it_16_cnu_37_in_1, msg_to_check_it_16_cnu_37_in_2, msg_to_check_it_16_cnu_37_in_3, msg_to_check_it_16_cnu_37_in_4, msg_to_check_it_16_cnu_37_in_5, msg_to_check_it_16_cnu_38_in_0, msg_to_check_it_16_cnu_38_in_1, msg_to_check_it_16_cnu_38_in_2, msg_to_check_it_16_cnu_38_in_3, msg_to_check_it_16_cnu_38_in_4, msg_to_check_it_16_cnu_38_in_5, msg_to_check_it_16_cnu_39_in_0, msg_to_check_it_16_cnu_39_in_1, msg_to_check_it_16_cnu_39_in_2, msg_to_check_it_16_cnu_39_in_3, msg_to_check_it_16_cnu_39_in_4, msg_to_check_it_16_cnu_39_in_5, msg_to_check_it_16_cnu_40_in_0, msg_to_check_it_16_cnu_40_in_1, msg_to_check_it_16_cnu_40_in_2, msg_to_check_it_16_cnu_40_in_3, msg_to_check_it_16_cnu_40_in_4, msg_to_check_it_16_cnu_40_in_5, msg_to_check_it_16_cnu_41_in_0, msg_to_check_it_16_cnu_41_in_1, msg_to_check_it_16_cnu_41_in_2, msg_to_check_it_16_cnu_41_in_3, msg_to_check_it_16_cnu_41_in_4, msg_to_check_it_16_cnu_41_in_5, msg_to_check_it_16_cnu_42_in_0, msg_to_check_it_16_cnu_42_in_1, msg_to_check_it_16_cnu_42_in_2, msg_to_check_it_16_cnu_42_in_3, msg_to_check_it_16_cnu_42_in_4, msg_to_check_it_16_cnu_42_in_5, msg_to_check_it_16_cnu_43_in_0, msg_to_check_it_16_cnu_43_in_1, msg_to_check_it_16_cnu_43_in_2, msg_to_check_it_16_cnu_43_in_3, msg_to_check_it_16_cnu_43_in_4, msg_to_check_it_16_cnu_43_in_5, msg_to_check_it_16_cnu_44_in_0, msg_to_check_it_16_cnu_44_in_1, msg_to_check_it_16_cnu_44_in_2, msg_to_check_it_16_cnu_44_in_3, msg_to_check_it_16_cnu_44_in_4, msg_to_check_it_16_cnu_44_in_5, msg_to_check_it_16_cnu_45_in_0, msg_to_check_it_16_cnu_45_in_1, msg_to_check_it_16_cnu_45_in_2, msg_to_check_it_16_cnu_45_in_3, msg_to_check_it_16_cnu_45_in_4, msg_to_check_it_16_cnu_45_in_5, msg_to_check_it_16_cnu_46_in_0, msg_to_check_it_16_cnu_46_in_1, msg_to_check_it_16_cnu_46_in_2, msg_to_check_it_16_cnu_46_in_3, msg_to_check_it_16_cnu_46_in_4, msg_to_check_it_16_cnu_46_in_5, msg_to_check_it_16_cnu_47_in_0, msg_to_check_it_16_cnu_47_in_1, msg_to_check_it_16_cnu_47_in_2, msg_to_check_it_16_cnu_47_in_3, msg_to_check_it_16_cnu_47_in_4, msg_to_check_it_16_cnu_47_in_5, msg_to_check_it_16_cnu_48_in_0, msg_to_check_it_16_cnu_48_in_1, msg_to_check_it_16_cnu_48_in_2, msg_to_check_it_16_cnu_48_in_3, msg_to_check_it_16_cnu_48_in_4, msg_to_check_it_16_cnu_48_in_5, msg_to_check_it_16_cnu_49_in_0, msg_to_check_it_16_cnu_49_in_1, msg_to_check_it_16_cnu_49_in_2, msg_to_check_it_16_cnu_49_in_3, msg_to_check_it_16_cnu_49_in_4, msg_to_check_it_16_cnu_49_in_5, msg_to_check_it_16_cnu_50_in_0, msg_to_check_it_16_cnu_50_in_1, msg_to_check_it_16_cnu_50_in_2, msg_to_check_it_16_cnu_50_in_3, msg_to_check_it_16_cnu_50_in_4, msg_to_check_it_16_cnu_50_in_5, msg_to_check_it_16_cnu_51_in_0, msg_to_check_it_16_cnu_51_in_1, msg_to_check_it_16_cnu_51_in_2, msg_to_check_it_16_cnu_51_in_3, msg_to_check_it_16_cnu_51_in_4, msg_to_check_it_16_cnu_51_in_5, msg_to_check_it_16_cnu_52_in_0, msg_to_check_it_16_cnu_52_in_1, msg_to_check_it_16_cnu_52_in_2, msg_to_check_it_16_cnu_52_in_3, msg_to_check_it_16_cnu_52_in_4, msg_to_check_it_16_cnu_52_in_5, msg_to_check_it_16_cnu_53_in_0, msg_to_check_it_16_cnu_53_in_1, msg_to_check_it_16_cnu_53_in_2, msg_to_check_it_16_cnu_53_in_3, msg_to_check_it_16_cnu_53_in_4, msg_to_check_it_16_cnu_53_in_5, msg_to_check_it_16_cnu_54_in_0, msg_to_check_it_16_cnu_54_in_1, msg_to_check_it_16_cnu_54_in_2, msg_to_check_it_16_cnu_54_in_3, msg_to_check_it_16_cnu_54_in_4, msg_to_check_it_16_cnu_54_in_5, msg_to_check_it_16_cnu_55_in_0, msg_to_check_it_16_cnu_55_in_1, msg_to_check_it_16_cnu_55_in_2, msg_to_check_it_16_cnu_55_in_3, msg_to_check_it_16_cnu_55_in_4, msg_to_check_it_16_cnu_55_in_5, msg_to_check_it_16_cnu_56_in_0, msg_to_check_it_16_cnu_56_in_1, msg_to_check_it_16_cnu_56_in_2, msg_to_check_it_16_cnu_56_in_3, msg_to_check_it_16_cnu_56_in_4, msg_to_check_it_16_cnu_56_in_5, msg_to_check_it_16_cnu_57_in_0, msg_to_check_it_16_cnu_57_in_1, msg_to_check_it_16_cnu_57_in_2, msg_to_check_it_16_cnu_57_in_3, msg_to_check_it_16_cnu_57_in_4, msg_to_check_it_16_cnu_57_in_5, msg_to_check_it_16_cnu_58_in_0, msg_to_check_it_16_cnu_58_in_1, msg_to_check_it_16_cnu_58_in_2, msg_to_check_it_16_cnu_58_in_3, msg_to_check_it_16_cnu_58_in_4, msg_to_check_it_16_cnu_58_in_5, msg_to_check_it_16_cnu_59_in_0, msg_to_check_it_16_cnu_59_in_1, msg_to_check_it_16_cnu_59_in_2, msg_to_check_it_16_cnu_59_in_3, msg_to_check_it_16_cnu_59_in_4, msg_to_check_it_16_cnu_59_in_5, msg_to_check_it_16_cnu_60_in_0, msg_to_check_it_16_cnu_60_in_1, msg_to_check_it_16_cnu_60_in_2, msg_to_check_it_16_cnu_60_in_3, msg_to_check_it_16_cnu_60_in_4, msg_to_check_it_16_cnu_60_in_5, msg_to_check_it_16_cnu_61_in_0, msg_to_check_it_16_cnu_61_in_1, msg_to_check_it_16_cnu_61_in_2, msg_to_check_it_16_cnu_61_in_3, msg_to_check_it_16_cnu_61_in_4, msg_to_check_it_16_cnu_61_in_5, msg_to_check_it_16_cnu_62_in_0, msg_to_check_it_16_cnu_62_in_1, msg_to_check_it_16_cnu_62_in_2, msg_to_check_it_16_cnu_62_in_3, msg_to_check_it_16_cnu_62_in_4, msg_to_check_it_16_cnu_62_in_5, msg_to_check_it_16_cnu_63_in_0, msg_to_check_it_16_cnu_63_in_1, msg_to_check_it_16_cnu_63_in_2, msg_to_check_it_16_cnu_63_in_3, msg_to_check_it_16_cnu_63_in_4, msg_to_check_it_16_cnu_63_in_5, msg_to_check_it_16_cnu_64_in_0, msg_to_check_it_16_cnu_64_in_1, msg_to_check_it_16_cnu_64_in_2, msg_to_check_it_16_cnu_64_in_3, msg_to_check_it_16_cnu_64_in_4, msg_to_check_it_16_cnu_64_in_5, msg_to_check_it_16_cnu_65_in_0, msg_to_check_it_16_cnu_65_in_1, msg_to_check_it_16_cnu_65_in_2, msg_to_check_it_16_cnu_65_in_3, msg_to_check_it_16_cnu_65_in_4, msg_to_check_it_16_cnu_65_in_5, msg_to_check_it_16_cnu_66_in_0, msg_to_check_it_16_cnu_66_in_1, msg_to_check_it_16_cnu_66_in_2, msg_to_check_it_16_cnu_66_in_3, msg_to_check_it_16_cnu_66_in_4, msg_to_check_it_16_cnu_66_in_5, msg_to_check_it_16_cnu_67_in_0, msg_to_check_it_16_cnu_67_in_1, msg_to_check_it_16_cnu_67_in_2, msg_to_check_it_16_cnu_67_in_3, msg_to_check_it_16_cnu_67_in_4, msg_to_check_it_16_cnu_67_in_5, msg_to_check_it_16_cnu_68_in_0, msg_to_check_it_16_cnu_68_in_1, msg_to_check_it_16_cnu_68_in_2, msg_to_check_it_16_cnu_68_in_3, msg_to_check_it_16_cnu_68_in_4, msg_to_check_it_16_cnu_68_in_5, msg_to_check_it_16_cnu_69_in_0, msg_to_check_it_16_cnu_69_in_1, msg_to_check_it_16_cnu_69_in_2, msg_to_check_it_16_cnu_69_in_3, msg_to_check_it_16_cnu_69_in_4, msg_to_check_it_16_cnu_69_in_5, msg_to_check_it_16_cnu_70_in_0, msg_to_check_it_16_cnu_70_in_1, msg_to_check_it_16_cnu_70_in_2, msg_to_check_it_16_cnu_70_in_3, msg_to_check_it_16_cnu_70_in_4, msg_to_check_it_16_cnu_70_in_5, msg_to_check_it_16_cnu_71_in_0, msg_to_check_it_16_cnu_71_in_1, msg_to_check_it_16_cnu_71_in_2, msg_to_check_it_16_cnu_71_in_3, msg_to_check_it_16_cnu_71_in_4, msg_to_check_it_16_cnu_71_in_5, msg_to_check_it_16_cnu_72_in_0, msg_to_check_it_16_cnu_72_in_1, msg_to_check_it_16_cnu_72_in_2, msg_to_check_it_16_cnu_72_in_3, msg_to_check_it_16_cnu_72_in_4, msg_to_check_it_16_cnu_72_in_5, msg_to_check_it_16_cnu_73_in_0, msg_to_check_it_16_cnu_73_in_1, msg_to_check_it_16_cnu_73_in_2, msg_to_check_it_16_cnu_73_in_3, msg_to_check_it_16_cnu_73_in_4, msg_to_check_it_16_cnu_73_in_5, msg_to_check_it_16_cnu_74_in_0, msg_to_check_it_16_cnu_74_in_1, msg_to_check_it_16_cnu_74_in_2, msg_to_check_it_16_cnu_74_in_3, msg_to_check_it_16_cnu_74_in_4, msg_to_check_it_16_cnu_74_in_5, msg_to_check_it_16_cnu_75_in_0, msg_to_check_it_16_cnu_75_in_1, msg_to_check_it_16_cnu_75_in_2, msg_to_check_it_16_cnu_75_in_3, msg_to_check_it_16_cnu_75_in_4, msg_to_check_it_16_cnu_75_in_5, msg_to_check_it_16_cnu_76_in_0, msg_to_check_it_16_cnu_76_in_1, msg_to_check_it_16_cnu_76_in_2, msg_to_check_it_16_cnu_76_in_3, msg_to_check_it_16_cnu_76_in_4, msg_to_check_it_16_cnu_76_in_5, msg_to_check_it_16_cnu_77_in_0, msg_to_check_it_16_cnu_77_in_1, msg_to_check_it_16_cnu_77_in_2, msg_to_check_it_16_cnu_77_in_3, msg_to_check_it_16_cnu_77_in_4, msg_to_check_it_16_cnu_77_in_5, msg_to_check_it_16_cnu_78_in_0, msg_to_check_it_16_cnu_78_in_1, msg_to_check_it_16_cnu_78_in_2, msg_to_check_it_16_cnu_78_in_3, msg_to_check_it_16_cnu_78_in_4, msg_to_check_it_16_cnu_78_in_5, msg_to_check_it_16_cnu_79_in_0, msg_to_check_it_16_cnu_79_in_1, msg_to_check_it_16_cnu_79_in_2, msg_to_check_it_16_cnu_79_in_3, msg_to_check_it_16_cnu_79_in_4, msg_to_check_it_16_cnu_79_in_5, msg_to_check_it_16_cnu_80_in_0, msg_to_check_it_16_cnu_80_in_1, msg_to_check_it_16_cnu_80_in_2, msg_to_check_it_16_cnu_80_in_3, msg_to_check_it_16_cnu_80_in_4, msg_to_check_it_16_cnu_80_in_5, msg_to_check_it_16_cnu_81_in_0, msg_to_check_it_16_cnu_81_in_1, msg_to_check_it_16_cnu_81_in_2, msg_to_check_it_16_cnu_81_in_3, msg_to_check_it_16_cnu_81_in_4, msg_to_check_it_16_cnu_81_in_5, msg_to_check_it_16_cnu_82_in_0, msg_to_check_it_16_cnu_82_in_1, msg_to_check_it_16_cnu_82_in_2, msg_to_check_it_16_cnu_82_in_3, msg_to_check_it_16_cnu_82_in_4, msg_to_check_it_16_cnu_82_in_5, msg_to_check_it_16_cnu_83_in_0, msg_to_check_it_16_cnu_83_in_1, msg_to_check_it_16_cnu_83_in_2, msg_to_check_it_16_cnu_83_in_3, msg_to_check_it_16_cnu_83_in_4, msg_to_check_it_16_cnu_83_in_5, msg_to_check_it_16_cnu_84_in_0, msg_to_check_it_16_cnu_84_in_1, msg_to_check_it_16_cnu_84_in_2, msg_to_check_it_16_cnu_84_in_3, msg_to_check_it_16_cnu_84_in_4, msg_to_check_it_16_cnu_84_in_5, msg_to_check_it_16_cnu_85_in_0, msg_to_check_it_16_cnu_85_in_1, msg_to_check_it_16_cnu_85_in_2, msg_to_check_it_16_cnu_85_in_3, msg_to_check_it_16_cnu_85_in_4, msg_to_check_it_16_cnu_85_in_5, msg_to_check_it_16_cnu_86_in_0, msg_to_check_it_16_cnu_86_in_1, msg_to_check_it_16_cnu_86_in_2, msg_to_check_it_16_cnu_86_in_3, msg_to_check_it_16_cnu_86_in_4, msg_to_check_it_16_cnu_86_in_5, msg_to_check_it_16_cnu_87_in_0, msg_to_check_it_16_cnu_87_in_1, msg_to_check_it_16_cnu_87_in_2, msg_to_check_it_16_cnu_87_in_3, msg_to_check_it_16_cnu_87_in_4, msg_to_check_it_16_cnu_87_in_5, msg_to_check_it_16_cnu_88_in_0, msg_to_check_it_16_cnu_88_in_1, msg_to_check_it_16_cnu_88_in_2, msg_to_check_it_16_cnu_88_in_3, msg_to_check_it_16_cnu_88_in_4, msg_to_check_it_16_cnu_88_in_5, msg_to_check_it_16_cnu_89_in_0, msg_to_check_it_16_cnu_89_in_1, msg_to_check_it_16_cnu_89_in_2, msg_to_check_it_16_cnu_89_in_3, msg_to_check_it_16_cnu_89_in_4, msg_to_check_it_16_cnu_89_in_5, msg_to_check_it_16_cnu_90_in_0, msg_to_check_it_16_cnu_90_in_1, msg_to_check_it_16_cnu_90_in_2, msg_to_check_it_16_cnu_90_in_3, msg_to_check_it_16_cnu_90_in_4, msg_to_check_it_16_cnu_90_in_5, msg_to_check_it_16_cnu_91_in_0, msg_to_check_it_16_cnu_91_in_1, msg_to_check_it_16_cnu_91_in_2, msg_to_check_it_16_cnu_91_in_3, msg_to_check_it_16_cnu_91_in_4, msg_to_check_it_16_cnu_91_in_5, msg_to_check_it_16_cnu_92_in_0, msg_to_check_it_16_cnu_92_in_1, msg_to_check_it_16_cnu_92_in_2, msg_to_check_it_16_cnu_92_in_3, msg_to_check_it_16_cnu_92_in_4, msg_to_check_it_16_cnu_92_in_5, msg_to_check_it_16_cnu_93_in_0, msg_to_check_it_16_cnu_93_in_1, msg_to_check_it_16_cnu_93_in_2, msg_to_check_it_16_cnu_93_in_3, msg_to_check_it_16_cnu_93_in_4, msg_to_check_it_16_cnu_93_in_5, msg_to_check_it_16_cnu_94_in_0, msg_to_check_it_16_cnu_94_in_1, msg_to_check_it_16_cnu_94_in_2, msg_to_check_it_16_cnu_94_in_3, msg_to_check_it_16_cnu_94_in_4, msg_to_check_it_16_cnu_94_in_5, msg_to_check_it_16_cnu_95_in_0, msg_to_check_it_16_cnu_95_in_1, msg_to_check_it_16_cnu_95_in_2, msg_to_check_it_16_cnu_95_in_3, msg_to_check_it_16_cnu_95_in_4, msg_to_check_it_16_cnu_95_in_5, msg_to_check_it_16_cnu_96_in_0, msg_to_check_it_16_cnu_96_in_1, msg_to_check_it_16_cnu_96_in_2, msg_to_check_it_16_cnu_96_in_3, msg_to_check_it_16_cnu_96_in_4, msg_to_check_it_16_cnu_96_in_5, msg_to_check_it_16_cnu_97_in_0, msg_to_check_it_16_cnu_97_in_1, msg_to_check_it_16_cnu_97_in_2, msg_to_check_it_16_cnu_97_in_3, msg_to_check_it_16_cnu_97_in_4, msg_to_check_it_16_cnu_97_in_5, msg_to_check_it_16_cnu_98_in_0, msg_to_check_it_16_cnu_98_in_1, msg_to_check_it_16_cnu_98_in_2, msg_to_check_it_16_cnu_98_in_3, msg_to_check_it_16_cnu_98_in_4, msg_to_check_it_16_cnu_98_in_5, msg_to_check_it_17_cnu_0_in_0, msg_to_check_it_17_cnu_0_in_1, msg_to_check_it_17_cnu_0_in_2, msg_to_check_it_17_cnu_0_in_3, msg_to_check_it_17_cnu_0_in_4, msg_to_check_it_17_cnu_0_in_5, msg_to_check_it_17_cnu_1_in_0, msg_to_check_it_17_cnu_1_in_1, msg_to_check_it_17_cnu_1_in_2, msg_to_check_it_17_cnu_1_in_3, msg_to_check_it_17_cnu_1_in_4, msg_to_check_it_17_cnu_1_in_5, msg_to_check_it_17_cnu_2_in_0, msg_to_check_it_17_cnu_2_in_1, msg_to_check_it_17_cnu_2_in_2, msg_to_check_it_17_cnu_2_in_3, msg_to_check_it_17_cnu_2_in_4, msg_to_check_it_17_cnu_2_in_5, msg_to_check_it_17_cnu_3_in_0, msg_to_check_it_17_cnu_3_in_1, msg_to_check_it_17_cnu_3_in_2, msg_to_check_it_17_cnu_3_in_3, msg_to_check_it_17_cnu_3_in_4, msg_to_check_it_17_cnu_3_in_5, msg_to_check_it_17_cnu_4_in_0, msg_to_check_it_17_cnu_4_in_1, msg_to_check_it_17_cnu_4_in_2, msg_to_check_it_17_cnu_4_in_3, msg_to_check_it_17_cnu_4_in_4, msg_to_check_it_17_cnu_4_in_5, msg_to_check_it_17_cnu_5_in_0, msg_to_check_it_17_cnu_5_in_1, msg_to_check_it_17_cnu_5_in_2, msg_to_check_it_17_cnu_5_in_3, msg_to_check_it_17_cnu_5_in_4, msg_to_check_it_17_cnu_5_in_5, msg_to_check_it_17_cnu_6_in_0, msg_to_check_it_17_cnu_6_in_1, msg_to_check_it_17_cnu_6_in_2, msg_to_check_it_17_cnu_6_in_3, msg_to_check_it_17_cnu_6_in_4, msg_to_check_it_17_cnu_6_in_5, msg_to_check_it_17_cnu_7_in_0, msg_to_check_it_17_cnu_7_in_1, msg_to_check_it_17_cnu_7_in_2, msg_to_check_it_17_cnu_7_in_3, msg_to_check_it_17_cnu_7_in_4, msg_to_check_it_17_cnu_7_in_5, msg_to_check_it_17_cnu_8_in_0, msg_to_check_it_17_cnu_8_in_1, msg_to_check_it_17_cnu_8_in_2, msg_to_check_it_17_cnu_8_in_3, msg_to_check_it_17_cnu_8_in_4, msg_to_check_it_17_cnu_8_in_5, msg_to_check_it_17_cnu_9_in_0, msg_to_check_it_17_cnu_9_in_1, msg_to_check_it_17_cnu_9_in_2, msg_to_check_it_17_cnu_9_in_3, msg_to_check_it_17_cnu_9_in_4, msg_to_check_it_17_cnu_9_in_5, msg_to_check_it_17_cnu_10_in_0, msg_to_check_it_17_cnu_10_in_1, msg_to_check_it_17_cnu_10_in_2, msg_to_check_it_17_cnu_10_in_3, msg_to_check_it_17_cnu_10_in_4, msg_to_check_it_17_cnu_10_in_5, msg_to_check_it_17_cnu_11_in_0, msg_to_check_it_17_cnu_11_in_1, msg_to_check_it_17_cnu_11_in_2, msg_to_check_it_17_cnu_11_in_3, msg_to_check_it_17_cnu_11_in_4, msg_to_check_it_17_cnu_11_in_5, msg_to_check_it_17_cnu_12_in_0, msg_to_check_it_17_cnu_12_in_1, msg_to_check_it_17_cnu_12_in_2, msg_to_check_it_17_cnu_12_in_3, msg_to_check_it_17_cnu_12_in_4, msg_to_check_it_17_cnu_12_in_5, msg_to_check_it_17_cnu_13_in_0, msg_to_check_it_17_cnu_13_in_1, msg_to_check_it_17_cnu_13_in_2, msg_to_check_it_17_cnu_13_in_3, msg_to_check_it_17_cnu_13_in_4, msg_to_check_it_17_cnu_13_in_5, msg_to_check_it_17_cnu_14_in_0, msg_to_check_it_17_cnu_14_in_1, msg_to_check_it_17_cnu_14_in_2, msg_to_check_it_17_cnu_14_in_3, msg_to_check_it_17_cnu_14_in_4, msg_to_check_it_17_cnu_14_in_5, msg_to_check_it_17_cnu_15_in_0, msg_to_check_it_17_cnu_15_in_1, msg_to_check_it_17_cnu_15_in_2, msg_to_check_it_17_cnu_15_in_3, msg_to_check_it_17_cnu_15_in_4, msg_to_check_it_17_cnu_15_in_5, msg_to_check_it_17_cnu_16_in_0, msg_to_check_it_17_cnu_16_in_1, msg_to_check_it_17_cnu_16_in_2, msg_to_check_it_17_cnu_16_in_3, msg_to_check_it_17_cnu_16_in_4, msg_to_check_it_17_cnu_16_in_5, msg_to_check_it_17_cnu_17_in_0, msg_to_check_it_17_cnu_17_in_1, msg_to_check_it_17_cnu_17_in_2, msg_to_check_it_17_cnu_17_in_3, msg_to_check_it_17_cnu_17_in_4, msg_to_check_it_17_cnu_17_in_5, msg_to_check_it_17_cnu_18_in_0, msg_to_check_it_17_cnu_18_in_1, msg_to_check_it_17_cnu_18_in_2, msg_to_check_it_17_cnu_18_in_3, msg_to_check_it_17_cnu_18_in_4, msg_to_check_it_17_cnu_18_in_5, msg_to_check_it_17_cnu_19_in_0, msg_to_check_it_17_cnu_19_in_1, msg_to_check_it_17_cnu_19_in_2, msg_to_check_it_17_cnu_19_in_3, msg_to_check_it_17_cnu_19_in_4, msg_to_check_it_17_cnu_19_in_5, msg_to_check_it_17_cnu_20_in_0, msg_to_check_it_17_cnu_20_in_1, msg_to_check_it_17_cnu_20_in_2, msg_to_check_it_17_cnu_20_in_3, msg_to_check_it_17_cnu_20_in_4, msg_to_check_it_17_cnu_20_in_5, msg_to_check_it_17_cnu_21_in_0, msg_to_check_it_17_cnu_21_in_1, msg_to_check_it_17_cnu_21_in_2, msg_to_check_it_17_cnu_21_in_3, msg_to_check_it_17_cnu_21_in_4, msg_to_check_it_17_cnu_21_in_5, msg_to_check_it_17_cnu_22_in_0, msg_to_check_it_17_cnu_22_in_1, msg_to_check_it_17_cnu_22_in_2, msg_to_check_it_17_cnu_22_in_3, msg_to_check_it_17_cnu_22_in_4, msg_to_check_it_17_cnu_22_in_5, msg_to_check_it_17_cnu_23_in_0, msg_to_check_it_17_cnu_23_in_1, msg_to_check_it_17_cnu_23_in_2, msg_to_check_it_17_cnu_23_in_3, msg_to_check_it_17_cnu_23_in_4, msg_to_check_it_17_cnu_23_in_5, msg_to_check_it_17_cnu_24_in_0, msg_to_check_it_17_cnu_24_in_1, msg_to_check_it_17_cnu_24_in_2, msg_to_check_it_17_cnu_24_in_3, msg_to_check_it_17_cnu_24_in_4, msg_to_check_it_17_cnu_24_in_5, msg_to_check_it_17_cnu_25_in_0, msg_to_check_it_17_cnu_25_in_1, msg_to_check_it_17_cnu_25_in_2, msg_to_check_it_17_cnu_25_in_3, msg_to_check_it_17_cnu_25_in_4, msg_to_check_it_17_cnu_25_in_5, msg_to_check_it_17_cnu_26_in_0, msg_to_check_it_17_cnu_26_in_1, msg_to_check_it_17_cnu_26_in_2, msg_to_check_it_17_cnu_26_in_3, msg_to_check_it_17_cnu_26_in_4, msg_to_check_it_17_cnu_26_in_5, msg_to_check_it_17_cnu_27_in_0, msg_to_check_it_17_cnu_27_in_1, msg_to_check_it_17_cnu_27_in_2, msg_to_check_it_17_cnu_27_in_3, msg_to_check_it_17_cnu_27_in_4, msg_to_check_it_17_cnu_27_in_5, msg_to_check_it_17_cnu_28_in_0, msg_to_check_it_17_cnu_28_in_1, msg_to_check_it_17_cnu_28_in_2, msg_to_check_it_17_cnu_28_in_3, msg_to_check_it_17_cnu_28_in_4, msg_to_check_it_17_cnu_28_in_5, msg_to_check_it_17_cnu_29_in_0, msg_to_check_it_17_cnu_29_in_1, msg_to_check_it_17_cnu_29_in_2, msg_to_check_it_17_cnu_29_in_3, msg_to_check_it_17_cnu_29_in_4, msg_to_check_it_17_cnu_29_in_5, msg_to_check_it_17_cnu_30_in_0, msg_to_check_it_17_cnu_30_in_1, msg_to_check_it_17_cnu_30_in_2, msg_to_check_it_17_cnu_30_in_3, msg_to_check_it_17_cnu_30_in_4, msg_to_check_it_17_cnu_30_in_5, msg_to_check_it_17_cnu_31_in_0, msg_to_check_it_17_cnu_31_in_1, msg_to_check_it_17_cnu_31_in_2, msg_to_check_it_17_cnu_31_in_3, msg_to_check_it_17_cnu_31_in_4, msg_to_check_it_17_cnu_31_in_5, msg_to_check_it_17_cnu_32_in_0, msg_to_check_it_17_cnu_32_in_1, msg_to_check_it_17_cnu_32_in_2, msg_to_check_it_17_cnu_32_in_3, msg_to_check_it_17_cnu_32_in_4, msg_to_check_it_17_cnu_32_in_5, msg_to_check_it_17_cnu_33_in_0, msg_to_check_it_17_cnu_33_in_1, msg_to_check_it_17_cnu_33_in_2, msg_to_check_it_17_cnu_33_in_3, msg_to_check_it_17_cnu_33_in_4, msg_to_check_it_17_cnu_33_in_5, msg_to_check_it_17_cnu_34_in_0, msg_to_check_it_17_cnu_34_in_1, msg_to_check_it_17_cnu_34_in_2, msg_to_check_it_17_cnu_34_in_3, msg_to_check_it_17_cnu_34_in_4, msg_to_check_it_17_cnu_34_in_5, msg_to_check_it_17_cnu_35_in_0, msg_to_check_it_17_cnu_35_in_1, msg_to_check_it_17_cnu_35_in_2, msg_to_check_it_17_cnu_35_in_3, msg_to_check_it_17_cnu_35_in_4, msg_to_check_it_17_cnu_35_in_5, msg_to_check_it_17_cnu_36_in_0, msg_to_check_it_17_cnu_36_in_1, msg_to_check_it_17_cnu_36_in_2, msg_to_check_it_17_cnu_36_in_3, msg_to_check_it_17_cnu_36_in_4, msg_to_check_it_17_cnu_36_in_5, msg_to_check_it_17_cnu_37_in_0, msg_to_check_it_17_cnu_37_in_1, msg_to_check_it_17_cnu_37_in_2, msg_to_check_it_17_cnu_37_in_3, msg_to_check_it_17_cnu_37_in_4, msg_to_check_it_17_cnu_37_in_5, msg_to_check_it_17_cnu_38_in_0, msg_to_check_it_17_cnu_38_in_1, msg_to_check_it_17_cnu_38_in_2, msg_to_check_it_17_cnu_38_in_3, msg_to_check_it_17_cnu_38_in_4, msg_to_check_it_17_cnu_38_in_5, msg_to_check_it_17_cnu_39_in_0, msg_to_check_it_17_cnu_39_in_1, msg_to_check_it_17_cnu_39_in_2, msg_to_check_it_17_cnu_39_in_3, msg_to_check_it_17_cnu_39_in_4, msg_to_check_it_17_cnu_39_in_5, msg_to_check_it_17_cnu_40_in_0, msg_to_check_it_17_cnu_40_in_1, msg_to_check_it_17_cnu_40_in_2, msg_to_check_it_17_cnu_40_in_3, msg_to_check_it_17_cnu_40_in_4, msg_to_check_it_17_cnu_40_in_5, msg_to_check_it_17_cnu_41_in_0, msg_to_check_it_17_cnu_41_in_1, msg_to_check_it_17_cnu_41_in_2, msg_to_check_it_17_cnu_41_in_3, msg_to_check_it_17_cnu_41_in_4, msg_to_check_it_17_cnu_41_in_5, msg_to_check_it_17_cnu_42_in_0, msg_to_check_it_17_cnu_42_in_1, msg_to_check_it_17_cnu_42_in_2, msg_to_check_it_17_cnu_42_in_3, msg_to_check_it_17_cnu_42_in_4, msg_to_check_it_17_cnu_42_in_5, msg_to_check_it_17_cnu_43_in_0, msg_to_check_it_17_cnu_43_in_1, msg_to_check_it_17_cnu_43_in_2, msg_to_check_it_17_cnu_43_in_3, msg_to_check_it_17_cnu_43_in_4, msg_to_check_it_17_cnu_43_in_5, msg_to_check_it_17_cnu_44_in_0, msg_to_check_it_17_cnu_44_in_1, msg_to_check_it_17_cnu_44_in_2, msg_to_check_it_17_cnu_44_in_3, msg_to_check_it_17_cnu_44_in_4, msg_to_check_it_17_cnu_44_in_5, msg_to_check_it_17_cnu_45_in_0, msg_to_check_it_17_cnu_45_in_1, msg_to_check_it_17_cnu_45_in_2, msg_to_check_it_17_cnu_45_in_3, msg_to_check_it_17_cnu_45_in_4, msg_to_check_it_17_cnu_45_in_5, msg_to_check_it_17_cnu_46_in_0, msg_to_check_it_17_cnu_46_in_1, msg_to_check_it_17_cnu_46_in_2, msg_to_check_it_17_cnu_46_in_3, msg_to_check_it_17_cnu_46_in_4, msg_to_check_it_17_cnu_46_in_5, msg_to_check_it_17_cnu_47_in_0, msg_to_check_it_17_cnu_47_in_1, msg_to_check_it_17_cnu_47_in_2, msg_to_check_it_17_cnu_47_in_3, msg_to_check_it_17_cnu_47_in_4, msg_to_check_it_17_cnu_47_in_5, msg_to_check_it_17_cnu_48_in_0, msg_to_check_it_17_cnu_48_in_1, msg_to_check_it_17_cnu_48_in_2, msg_to_check_it_17_cnu_48_in_3, msg_to_check_it_17_cnu_48_in_4, msg_to_check_it_17_cnu_48_in_5, msg_to_check_it_17_cnu_49_in_0, msg_to_check_it_17_cnu_49_in_1, msg_to_check_it_17_cnu_49_in_2, msg_to_check_it_17_cnu_49_in_3, msg_to_check_it_17_cnu_49_in_4, msg_to_check_it_17_cnu_49_in_5, msg_to_check_it_17_cnu_50_in_0, msg_to_check_it_17_cnu_50_in_1, msg_to_check_it_17_cnu_50_in_2, msg_to_check_it_17_cnu_50_in_3, msg_to_check_it_17_cnu_50_in_4, msg_to_check_it_17_cnu_50_in_5, msg_to_check_it_17_cnu_51_in_0, msg_to_check_it_17_cnu_51_in_1, msg_to_check_it_17_cnu_51_in_2, msg_to_check_it_17_cnu_51_in_3, msg_to_check_it_17_cnu_51_in_4, msg_to_check_it_17_cnu_51_in_5, msg_to_check_it_17_cnu_52_in_0, msg_to_check_it_17_cnu_52_in_1, msg_to_check_it_17_cnu_52_in_2, msg_to_check_it_17_cnu_52_in_3, msg_to_check_it_17_cnu_52_in_4, msg_to_check_it_17_cnu_52_in_5, msg_to_check_it_17_cnu_53_in_0, msg_to_check_it_17_cnu_53_in_1, msg_to_check_it_17_cnu_53_in_2, msg_to_check_it_17_cnu_53_in_3, msg_to_check_it_17_cnu_53_in_4, msg_to_check_it_17_cnu_53_in_5, msg_to_check_it_17_cnu_54_in_0, msg_to_check_it_17_cnu_54_in_1, msg_to_check_it_17_cnu_54_in_2, msg_to_check_it_17_cnu_54_in_3, msg_to_check_it_17_cnu_54_in_4, msg_to_check_it_17_cnu_54_in_5, msg_to_check_it_17_cnu_55_in_0, msg_to_check_it_17_cnu_55_in_1, msg_to_check_it_17_cnu_55_in_2, msg_to_check_it_17_cnu_55_in_3, msg_to_check_it_17_cnu_55_in_4, msg_to_check_it_17_cnu_55_in_5, msg_to_check_it_17_cnu_56_in_0, msg_to_check_it_17_cnu_56_in_1, msg_to_check_it_17_cnu_56_in_2, msg_to_check_it_17_cnu_56_in_3, msg_to_check_it_17_cnu_56_in_4, msg_to_check_it_17_cnu_56_in_5, msg_to_check_it_17_cnu_57_in_0, msg_to_check_it_17_cnu_57_in_1, msg_to_check_it_17_cnu_57_in_2, msg_to_check_it_17_cnu_57_in_3, msg_to_check_it_17_cnu_57_in_4, msg_to_check_it_17_cnu_57_in_5, msg_to_check_it_17_cnu_58_in_0, msg_to_check_it_17_cnu_58_in_1, msg_to_check_it_17_cnu_58_in_2, msg_to_check_it_17_cnu_58_in_3, msg_to_check_it_17_cnu_58_in_4, msg_to_check_it_17_cnu_58_in_5, msg_to_check_it_17_cnu_59_in_0, msg_to_check_it_17_cnu_59_in_1, msg_to_check_it_17_cnu_59_in_2, msg_to_check_it_17_cnu_59_in_3, msg_to_check_it_17_cnu_59_in_4, msg_to_check_it_17_cnu_59_in_5, msg_to_check_it_17_cnu_60_in_0, msg_to_check_it_17_cnu_60_in_1, msg_to_check_it_17_cnu_60_in_2, msg_to_check_it_17_cnu_60_in_3, msg_to_check_it_17_cnu_60_in_4, msg_to_check_it_17_cnu_60_in_5, msg_to_check_it_17_cnu_61_in_0, msg_to_check_it_17_cnu_61_in_1, msg_to_check_it_17_cnu_61_in_2, msg_to_check_it_17_cnu_61_in_3, msg_to_check_it_17_cnu_61_in_4, msg_to_check_it_17_cnu_61_in_5, msg_to_check_it_17_cnu_62_in_0, msg_to_check_it_17_cnu_62_in_1, msg_to_check_it_17_cnu_62_in_2, msg_to_check_it_17_cnu_62_in_3, msg_to_check_it_17_cnu_62_in_4, msg_to_check_it_17_cnu_62_in_5, msg_to_check_it_17_cnu_63_in_0, msg_to_check_it_17_cnu_63_in_1, msg_to_check_it_17_cnu_63_in_2, msg_to_check_it_17_cnu_63_in_3, msg_to_check_it_17_cnu_63_in_4, msg_to_check_it_17_cnu_63_in_5, msg_to_check_it_17_cnu_64_in_0, msg_to_check_it_17_cnu_64_in_1, msg_to_check_it_17_cnu_64_in_2, msg_to_check_it_17_cnu_64_in_3, msg_to_check_it_17_cnu_64_in_4, msg_to_check_it_17_cnu_64_in_5, msg_to_check_it_17_cnu_65_in_0, msg_to_check_it_17_cnu_65_in_1, msg_to_check_it_17_cnu_65_in_2, msg_to_check_it_17_cnu_65_in_3, msg_to_check_it_17_cnu_65_in_4, msg_to_check_it_17_cnu_65_in_5, msg_to_check_it_17_cnu_66_in_0, msg_to_check_it_17_cnu_66_in_1, msg_to_check_it_17_cnu_66_in_2, msg_to_check_it_17_cnu_66_in_3, msg_to_check_it_17_cnu_66_in_4, msg_to_check_it_17_cnu_66_in_5, msg_to_check_it_17_cnu_67_in_0, msg_to_check_it_17_cnu_67_in_1, msg_to_check_it_17_cnu_67_in_2, msg_to_check_it_17_cnu_67_in_3, msg_to_check_it_17_cnu_67_in_4, msg_to_check_it_17_cnu_67_in_5, msg_to_check_it_17_cnu_68_in_0, msg_to_check_it_17_cnu_68_in_1, msg_to_check_it_17_cnu_68_in_2, msg_to_check_it_17_cnu_68_in_3, msg_to_check_it_17_cnu_68_in_4, msg_to_check_it_17_cnu_68_in_5, msg_to_check_it_17_cnu_69_in_0, msg_to_check_it_17_cnu_69_in_1, msg_to_check_it_17_cnu_69_in_2, msg_to_check_it_17_cnu_69_in_3, msg_to_check_it_17_cnu_69_in_4, msg_to_check_it_17_cnu_69_in_5, msg_to_check_it_17_cnu_70_in_0, msg_to_check_it_17_cnu_70_in_1, msg_to_check_it_17_cnu_70_in_2, msg_to_check_it_17_cnu_70_in_3, msg_to_check_it_17_cnu_70_in_4, msg_to_check_it_17_cnu_70_in_5, msg_to_check_it_17_cnu_71_in_0, msg_to_check_it_17_cnu_71_in_1, msg_to_check_it_17_cnu_71_in_2, msg_to_check_it_17_cnu_71_in_3, msg_to_check_it_17_cnu_71_in_4, msg_to_check_it_17_cnu_71_in_5, msg_to_check_it_17_cnu_72_in_0, msg_to_check_it_17_cnu_72_in_1, msg_to_check_it_17_cnu_72_in_2, msg_to_check_it_17_cnu_72_in_3, msg_to_check_it_17_cnu_72_in_4, msg_to_check_it_17_cnu_72_in_5, msg_to_check_it_17_cnu_73_in_0, msg_to_check_it_17_cnu_73_in_1, msg_to_check_it_17_cnu_73_in_2, msg_to_check_it_17_cnu_73_in_3, msg_to_check_it_17_cnu_73_in_4, msg_to_check_it_17_cnu_73_in_5, msg_to_check_it_17_cnu_74_in_0, msg_to_check_it_17_cnu_74_in_1, msg_to_check_it_17_cnu_74_in_2, msg_to_check_it_17_cnu_74_in_3, msg_to_check_it_17_cnu_74_in_4, msg_to_check_it_17_cnu_74_in_5, msg_to_check_it_17_cnu_75_in_0, msg_to_check_it_17_cnu_75_in_1, msg_to_check_it_17_cnu_75_in_2, msg_to_check_it_17_cnu_75_in_3, msg_to_check_it_17_cnu_75_in_4, msg_to_check_it_17_cnu_75_in_5, msg_to_check_it_17_cnu_76_in_0, msg_to_check_it_17_cnu_76_in_1, msg_to_check_it_17_cnu_76_in_2, msg_to_check_it_17_cnu_76_in_3, msg_to_check_it_17_cnu_76_in_4, msg_to_check_it_17_cnu_76_in_5, msg_to_check_it_17_cnu_77_in_0, msg_to_check_it_17_cnu_77_in_1, msg_to_check_it_17_cnu_77_in_2, msg_to_check_it_17_cnu_77_in_3, msg_to_check_it_17_cnu_77_in_4, msg_to_check_it_17_cnu_77_in_5, msg_to_check_it_17_cnu_78_in_0, msg_to_check_it_17_cnu_78_in_1, msg_to_check_it_17_cnu_78_in_2, msg_to_check_it_17_cnu_78_in_3, msg_to_check_it_17_cnu_78_in_4, msg_to_check_it_17_cnu_78_in_5, msg_to_check_it_17_cnu_79_in_0, msg_to_check_it_17_cnu_79_in_1, msg_to_check_it_17_cnu_79_in_2, msg_to_check_it_17_cnu_79_in_3, msg_to_check_it_17_cnu_79_in_4, msg_to_check_it_17_cnu_79_in_5, msg_to_check_it_17_cnu_80_in_0, msg_to_check_it_17_cnu_80_in_1, msg_to_check_it_17_cnu_80_in_2, msg_to_check_it_17_cnu_80_in_3, msg_to_check_it_17_cnu_80_in_4, msg_to_check_it_17_cnu_80_in_5, msg_to_check_it_17_cnu_81_in_0, msg_to_check_it_17_cnu_81_in_1, msg_to_check_it_17_cnu_81_in_2, msg_to_check_it_17_cnu_81_in_3, msg_to_check_it_17_cnu_81_in_4, msg_to_check_it_17_cnu_81_in_5, msg_to_check_it_17_cnu_82_in_0, msg_to_check_it_17_cnu_82_in_1, msg_to_check_it_17_cnu_82_in_2, msg_to_check_it_17_cnu_82_in_3, msg_to_check_it_17_cnu_82_in_4, msg_to_check_it_17_cnu_82_in_5, msg_to_check_it_17_cnu_83_in_0, msg_to_check_it_17_cnu_83_in_1, msg_to_check_it_17_cnu_83_in_2, msg_to_check_it_17_cnu_83_in_3, msg_to_check_it_17_cnu_83_in_4, msg_to_check_it_17_cnu_83_in_5, msg_to_check_it_17_cnu_84_in_0, msg_to_check_it_17_cnu_84_in_1, msg_to_check_it_17_cnu_84_in_2, msg_to_check_it_17_cnu_84_in_3, msg_to_check_it_17_cnu_84_in_4, msg_to_check_it_17_cnu_84_in_5, msg_to_check_it_17_cnu_85_in_0, msg_to_check_it_17_cnu_85_in_1, msg_to_check_it_17_cnu_85_in_2, msg_to_check_it_17_cnu_85_in_3, msg_to_check_it_17_cnu_85_in_4, msg_to_check_it_17_cnu_85_in_5, msg_to_check_it_17_cnu_86_in_0, msg_to_check_it_17_cnu_86_in_1, msg_to_check_it_17_cnu_86_in_2, msg_to_check_it_17_cnu_86_in_3, msg_to_check_it_17_cnu_86_in_4, msg_to_check_it_17_cnu_86_in_5, msg_to_check_it_17_cnu_87_in_0, msg_to_check_it_17_cnu_87_in_1, msg_to_check_it_17_cnu_87_in_2, msg_to_check_it_17_cnu_87_in_3, msg_to_check_it_17_cnu_87_in_4, msg_to_check_it_17_cnu_87_in_5, msg_to_check_it_17_cnu_88_in_0, msg_to_check_it_17_cnu_88_in_1, msg_to_check_it_17_cnu_88_in_2, msg_to_check_it_17_cnu_88_in_3, msg_to_check_it_17_cnu_88_in_4, msg_to_check_it_17_cnu_88_in_5, msg_to_check_it_17_cnu_89_in_0, msg_to_check_it_17_cnu_89_in_1, msg_to_check_it_17_cnu_89_in_2, msg_to_check_it_17_cnu_89_in_3, msg_to_check_it_17_cnu_89_in_4, msg_to_check_it_17_cnu_89_in_5, msg_to_check_it_17_cnu_90_in_0, msg_to_check_it_17_cnu_90_in_1, msg_to_check_it_17_cnu_90_in_2, msg_to_check_it_17_cnu_90_in_3, msg_to_check_it_17_cnu_90_in_4, msg_to_check_it_17_cnu_90_in_5, msg_to_check_it_17_cnu_91_in_0, msg_to_check_it_17_cnu_91_in_1, msg_to_check_it_17_cnu_91_in_2, msg_to_check_it_17_cnu_91_in_3, msg_to_check_it_17_cnu_91_in_4, msg_to_check_it_17_cnu_91_in_5, msg_to_check_it_17_cnu_92_in_0, msg_to_check_it_17_cnu_92_in_1, msg_to_check_it_17_cnu_92_in_2, msg_to_check_it_17_cnu_92_in_3, msg_to_check_it_17_cnu_92_in_4, msg_to_check_it_17_cnu_92_in_5, msg_to_check_it_17_cnu_93_in_0, msg_to_check_it_17_cnu_93_in_1, msg_to_check_it_17_cnu_93_in_2, msg_to_check_it_17_cnu_93_in_3, msg_to_check_it_17_cnu_93_in_4, msg_to_check_it_17_cnu_93_in_5, msg_to_check_it_17_cnu_94_in_0, msg_to_check_it_17_cnu_94_in_1, msg_to_check_it_17_cnu_94_in_2, msg_to_check_it_17_cnu_94_in_3, msg_to_check_it_17_cnu_94_in_4, msg_to_check_it_17_cnu_94_in_5, msg_to_check_it_17_cnu_95_in_0, msg_to_check_it_17_cnu_95_in_1, msg_to_check_it_17_cnu_95_in_2, msg_to_check_it_17_cnu_95_in_3, msg_to_check_it_17_cnu_95_in_4, msg_to_check_it_17_cnu_95_in_5, msg_to_check_it_17_cnu_96_in_0, msg_to_check_it_17_cnu_96_in_1, msg_to_check_it_17_cnu_96_in_2, msg_to_check_it_17_cnu_96_in_3, msg_to_check_it_17_cnu_96_in_4, msg_to_check_it_17_cnu_96_in_5, msg_to_check_it_17_cnu_97_in_0, msg_to_check_it_17_cnu_97_in_1, msg_to_check_it_17_cnu_97_in_2, msg_to_check_it_17_cnu_97_in_3, msg_to_check_it_17_cnu_97_in_4, msg_to_check_it_17_cnu_97_in_5, msg_to_check_it_17_cnu_98_in_0, msg_to_check_it_17_cnu_98_in_1, msg_to_check_it_17_cnu_98_in_2, msg_to_check_it_17_cnu_98_in_3, msg_to_check_it_17_cnu_98_in_4, msg_to_check_it_17_cnu_98_in_5, msg_to_check_it_18_cnu_0_in_0, msg_to_check_it_18_cnu_0_in_1, msg_to_check_it_18_cnu_0_in_2, msg_to_check_it_18_cnu_0_in_3, msg_to_check_it_18_cnu_0_in_4, msg_to_check_it_18_cnu_0_in_5, msg_to_check_it_18_cnu_1_in_0, msg_to_check_it_18_cnu_1_in_1, msg_to_check_it_18_cnu_1_in_2, msg_to_check_it_18_cnu_1_in_3, msg_to_check_it_18_cnu_1_in_4, msg_to_check_it_18_cnu_1_in_5, msg_to_check_it_18_cnu_2_in_0, msg_to_check_it_18_cnu_2_in_1, msg_to_check_it_18_cnu_2_in_2, msg_to_check_it_18_cnu_2_in_3, msg_to_check_it_18_cnu_2_in_4, msg_to_check_it_18_cnu_2_in_5, msg_to_check_it_18_cnu_3_in_0, msg_to_check_it_18_cnu_3_in_1, msg_to_check_it_18_cnu_3_in_2, msg_to_check_it_18_cnu_3_in_3, msg_to_check_it_18_cnu_3_in_4, msg_to_check_it_18_cnu_3_in_5, msg_to_check_it_18_cnu_4_in_0, msg_to_check_it_18_cnu_4_in_1, msg_to_check_it_18_cnu_4_in_2, msg_to_check_it_18_cnu_4_in_3, msg_to_check_it_18_cnu_4_in_4, msg_to_check_it_18_cnu_4_in_5, msg_to_check_it_18_cnu_5_in_0, msg_to_check_it_18_cnu_5_in_1, msg_to_check_it_18_cnu_5_in_2, msg_to_check_it_18_cnu_5_in_3, msg_to_check_it_18_cnu_5_in_4, msg_to_check_it_18_cnu_5_in_5, msg_to_check_it_18_cnu_6_in_0, msg_to_check_it_18_cnu_6_in_1, msg_to_check_it_18_cnu_6_in_2, msg_to_check_it_18_cnu_6_in_3, msg_to_check_it_18_cnu_6_in_4, msg_to_check_it_18_cnu_6_in_5, msg_to_check_it_18_cnu_7_in_0, msg_to_check_it_18_cnu_7_in_1, msg_to_check_it_18_cnu_7_in_2, msg_to_check_it_18_cnu_7_in_3, msg_to_check_it_18_cnu_7_in_4, msg_to_check_it_18_cnu_7_in_5, msg_to_check_it_18_cnu_8_in_0, msg_to_check_it_18_cnu_8_in_1, msg_to_check_it_18_cnu_8_in_2, msg_to_check_it_18_cnu_8_in_3, msg_to_check_it_18_cnu_8_in_4, msg_to_check_it_18_cnu_8_in_5, msg_to_check_it_18_cnu_9_in_0, msg_to_check_it_18_cnu_9_in_1, msg_to_check_it_18_cnu_9_in_2, msg_to_check_it_18_cnu_9_in_3, msg_to_check_it_18_cnu_9_in_4, msg_to_check_it_18_cnu_9_in_5, msg_to_check_it_18_cnu_10_in_0, msg_to_check_it_18_cnu_10_in_1, msg_to_check_it_18_cnu_10_in_2, msg_to_check_it_18_cnu_10_in_3, msg_to_check_it_18_cnu_10_in_4, msg_to_check_it_18_cnu_10_in_5, msg_to_check_it_18_cnu_11_in_0, msg_to_check_it_18_cnu_11_in_1, msg_to_check_it_18_cnu_11_in_2, msg_to_check_it_18_cnu_11_in_3, msg_to_check_it_18_cnu_11_in_4, msg_to_check_it_18_cnu_11_in_5, msg_to_check_it_18_cnu_12_in_0, msg_to_check_it_18_cnu_12_in_1, msg_to_check_it_18_cnu_12_in_2, msg_to_check_it_18_cnu_12_in_3, msg_to_check_it_18_cnu_12_in_4, msg_to_check_it_18_cnu_12_in_5, msg_to_check_it_18_cnu_13_in_0, msg_to_check_it_18_cnu_13_in_1, msg_to_check_it_18_cnu_13_in_2, msg_to_check_it_18_cnu_13_in_3, msg_to_check_it_18_cnu_13_in_4, msg_to_check_it_18_cnu_13_in_5, msg_to_check_it_18_cnu_14_in_0, msg_to_check_it_18_cnu_14_in_1, msg_to_check_it_18_cnu_14_in_2, msg_to_check_it_18_cnu_14_in_3, msg_to_check_it_18_cnu_14_in_4, msg_to_check_it_18_cnu_14_in_5, msg_to_check_it_18_cnu_15_in_0, msg_to_check_it_18_cnu_15_in_1, msg_to_check_it_18_cnu_15_in_2, msg_to_check_it_18_cnu_15_in_3, msg_to_check_it_18_cnu_15_in_4, msg_to_check_it_18_cnu_15_in_5, msg_to_check_it_18_cnu_16_in_0, msg_to_check_it_18_cnu_16_in_1, msg_to_check_it_18_cnu_16_in_2, msg_to_check_it_18_cnu_16_in_3, msg_to_check_it_18_cnu_16_in_4, msg_to_check_it_18_cnu_16_in_5, msg_to_check_it_18_cnu_17_in_0, msg_to_check_it_18_cnu_17_in_1, msg_to_check_it_18_cnu_17_in_2, msg_to_check_it_18_cnu_17_in_3, msg_to_check_it_18_cnu_17_in_4, msg_to_check_it_18_cnu_17_in_5, msg_to_check_it_18_cnu_18_in_0, msg_to_check_it_18_cnu_18_in_1, msg_to_check_it_18_cnu_18_in_2, msg_to_check_it_18_cnu_18_in_3, msg_to_check_it_18_cnu_18_in_4, msg_to_check_it_18_cnu_18_in_5, msg_to_check_it_18_cnu_19_in_0, msg_to_check_it_18_cnu_19_in_1, msg_to_check_it_18_cnu_19_in_2, msg_to_check_it_18_cnu_19_in_3, msg_to_check_it_18_cnu_19_in_4, msg_to_check_it_18_cnu_19_in_5, msg_to_check_it_18_cnu_20_in_0, msg_to_check_it_18_cnu_20_in_1, msg_to_check_it_18_cnu_20_in_2, msg_to_check_it_18_cnu_20_in_3, msg_to_check_it_18_cnu_20_in_4, msg_to_check_it_18_cnu_20_in_5, msg_to_check_it_18_cnu_21_in_0, msg_to_check_it_18_cnu_21_in_1, msg_to_check_it_18_cnu_21_in_2, msg_to_check_it_18_cnu_21_in_3, msg_to_check_it_18_cnu_21_in_4, msg_to_check_it_18_cnu_21_in_5, msg_to_check_it_18_cnu_22_in_0, msg_to_check_it_18_cnu_22_in_1, msg_to_check_it_18_cnu_22_in_2, msg_to_check_it_18_cnu_22_in_3, msg_to_check_it_18_cnu_22_in_4, msg_to_check_it_18_cnu_22_in_5, msg_to_check_it_18_cnu_23_in_0, msg_to_check_it_18_cnu_23_in_1, msg_to_check_it_18_cnu_23_in_2, msg_to_check_it_18_cnu_23_in_3, msg_to_check_it_18_cnu_23_in_4, msg_to_check_it_18_cnu_23_in_5, msg_to_check_it_18_cnu_24_in_0, msg_to_check_it_18_cnu_24_in_1, msg_to_check_it_18_cnu_24_in_2, msg_to_check_it_18_cnu_24_in_3, msg_to_check_it_18_cnu_24_in_4, msg_to_check_it_18_cnu_24_in_5, msg_to_check_it_18_cnu_25_in_0, msg_to_check_it_18_cnu_25_in_1, msg_to_check_it_18_cnu_25_in_2, msg_to_check_it_18_cnu_25_in_3, msg_to_check_it_18_cnu_25_in_4, msg_to_check_it_18_cnu_25_in_5, msg_to_check_it_18_cnu_26_in_0, msg_to_check_it_18_cnu_26_in_1, msg_to_check_it_18_cnu_26_in_2, msg_to_check_it_18_cnu_26_in_3, msg_to_check_it_18_cnu_26_in_4, msg_to_check_it_18_cnu_26_in_5, msg_to_check_it_18_cnu_27_in_0, msg_to_check_it_18_cnu_27_in_1, msg_to_check_it_18_cnu_27_in_2, msg_to_check_it_18_cnu_27_in_3, msg_to_check_it_18_cnu_27_in_4, msg_to_check_it_18_cnu_27_in_5, msg_to_check_it_18_cnu_28_in_0, msg_to_check_it_18_cnu_28_in_1, msg_to_check_it_18_cnu_28_in_2, msg_to_check_it_18_cnu_28_in_3, msg_to_check_it_18_cnu_28_in_4, msg_to_check_it_18_cnu_28_in_5, msg_to_check_it_18_cnu_29_in_0, msg_to_check_it_18_cnu_29_in_1, msg_to_check_it_18_cnu_29_in_2, msg_to_check_it_18_cnu_29_in_3, msg_to_check_it_18_cnu_29_in_4, msg_to_check_it_18_cnu_29_in_5, msg_to_check_it_18_cnu_30_in_0, msg_to_check_it_18_cnu_30_in_1, msg_to_check_it_18_cnu_30_in_2, msg_to_check_it_18_cnu_30_in_3, msg_to_check_it_18_cnu_30_in_4, msg_to_check_it_18_cnu_30_in_5, msg_to_check_it_18_cnu_31_in_0, msg_to_check_it_18_cnu_31_in_1, msg_to_check_it_18_cnu_31_in_2, msg_to_check_it_18_cnu_31_in_3, msg_to_check_it_18_cnu_31_in_4, msg_to_check_it_18_cnu_31_in_5, msg_to_check_it_18_cnu_32_in_0, msg_to_check_it_18_cnu_32_in_1, msg_to_check_it_18_cnu_32_in_2, msg_to_check_it_18_cnu_32_in_3, msg_to_check_it_18_cnu_32_in_4, msg_to_check_it_18_cnu_32_in_5, msg_to_check_it_18_cnu_33_in_0, msg_to_check_it_18_cnu_33_in_1, msg_to_check_it_18_cnu_33_in_2, msg_to_check_it_18_cnu_33_in_3, msg_to_check_it_18_cnu_33_in_4, msg_to_check_it_18_cnu_33_in_5, msg_to_check_it_18_cnu_34_in_0, msg_to_check_it_18_cnu_34_in_1, msg_to_check_it_18_cnu_34_in_2, msg_to_check_it_18_cnu_34_in_3, msg_to_check_it_18_cnu_34_in_4, msg_to_check_it_18_cnu_34_in_5, msg_to_check_it_18_cnu_35_in_0, msg_to_check_it_18_cnu_35_in_1, msg_to_check_it_18_cnu_35_in_2, msg_to_check_it_18_cnu_35_in_3, msg_to_check_it_18_cnu_35_in_4, msg_to_check_it_18_cnu_35_in_5, msg_to_check_it_18_cnu_36_in_0, msg_to_check_it_18_cnu_36_in_1, msg_to_check_it_18_cnu_36_in_2, msg_to_check_it_18_cnu_36_in_3, msg_to_check_it_18_cnu_36_in_4, msg_to_check_it_18_cnu_36_in_5, msg_to_check_it_18_cnu_37_in_0, msg_to_check_it_18_cnu_37_in_1, msg_to_check_it_18_cnu_37_in_2, msg_to_check_it_18_cnu_37_in_3, msg_to_check_it_18_cnu_37_in_4, msg_to_check_it_18_cnu_37_in_5, msg_to_check_it_18_cnu_38_in_0, msg_to_check_it_18_cnu_38_in_1, msg_to_check_it_18_cnu_38_in_2, msg_to_check_it_18_cnu_38_in_3, msg_to_check_it_18_cnu_38_in_4, msg_to_check_it_18_cnu_38_in_5, msg_to_check_it_18_cnu_39_in_0, msg_to_check_it_18_cnu_39_in_1, msg_to_check_it_18_cnu_39_in_2, msg_to_check_it_18_cnu_39_in_3, msg_to_check_it_18_cnu_39_in_4, msg_to_check_it_18_cnu_39_in_5, msg_to_check_it_18_cnu_40_in_0, msg_to_check_it_18_cnu_40_in_1, msg_to_check_it_18_cnu_40_in_2, msg_to_check_it_18_cnu_40_in_3, msg_to_check_it_18_cnu_40_in_4, msg_to_check_it_18_cnu_40_in_5, msg_to_check_it_18_cnu_41_in_0, msg_to_check_it_18_cnu_41_in_1, msg_to_check_it_18_cnu_41_in_2, msg_to_check_it_18_cnu_41_in_3, msg_to_check_it_18_cnu_41_in_4, msg_to_check_it_18_cnu_41_in_5, msg_to_check_it_18_cnu_42_in_0, msg_to_check_it_18_cnu_42_in_1, msg_to_check_it_18_cnu_42_in_2, msg_to_check_it_18_cnu_42_in_3, msg_to_check_it_18_cnu_42_in_4, msg_to_check_it_18_cnu_42_in_5, msg_to_check_it_18_cnu_43_in_0, msg_to_check_it_18_cnu_43_in_1, msg_to_check_it_18_cnu_43_in_2, msg_to_check_it_18_cnu_43_in_3, msg_to_check_it_18_cnu_43_in_4, msg_to_check_it_18_cnu_43_in_5, msg_to_check_it_18_cnu_44_in_0, msg_to_check_it_18_cnu_44_in_1, msg_to_check_it_18_cnu_44_in_2, msg_to_check_it_18_cnu_44_in_3, msg_to_check_it_18_cnu_44_in_4, msg_to_check_it_18_cnu_44_in_5, msg_to_check_it_18_cnu_45_in_0, msg_to_check_it_18_cnu_45_in_1, msg_to_check_it_18_cnu_45_in_2, msg_to_check_it_18_cnu_45_in_3, msg_to_check_it_18_cnu_45_in_4, msg_to_check_it_18_cnu_45_in_5, msg_to_check_it_18_cnu_46_in_0, msg_to_check_it_18_cnu_46_in_1, msg_to_check_it_18_cnu_46_in_2, msg_to_check_it_18_cnu_46_in_3, msg_to_check_it_18_cnu_46_in_4, msg_to_check_it_18_cnu_46_in_5, msg_to_check_it_18_cnu_47_in_0, msg_to_check_it_18_cnu_47_in_1, msg_to_check_it_18_cnu_47_in_2, msg_to_check_it_18_cnu_47_in_3, msg_to_check_it_18_cnu_47_in_4, msg_to_check_it_18_cnu_47_in_5, msg_to_check_it_18_cnu_48_in_0, msg_to_check_it_18_cnu_48_in_1, msg_to_check_it_18_cnu_48_in_2, msg_to_check_it_18_cnu_48_in_3, msg_to_check_it_18_cnu_48_in_4, msg_to_check_it_18_cnu_48_in_5, msg_to_check_it_18_cnu_49_in_0, msg_to_check_it_18_cnu_49_in_1, msg_to_check_it_18_cnu_49_in_2, msg_to_check_it_18_cnu_49_in_3, msg_to_check_it_18_cnu_49_in_4, msg_to_check_it_18_cnu_49_in_5, msg_to_check_it_18_cnu_50_in_0, msg_to_check_it_18_cnu_50_in_1, msg_to_check_it_18_cnu_50_in_2, msg_to_check_it_18_cnu_50_in_3, msg_to_check_it_18_cnu_50_in_4, msg_to_check_it_18_cnu_50_in_5, msg_to_check_it_18_cnu_51_in_0, msg_to_check_it_18_cnu_51_in_1, msg_to_check_it_18_cnu_51_in_2, msg_to_check_it_18_cnu_51_in_3, msg_to_check_it_18_cnu_51_in_4, msg_to_check_it_18_cnu_51_in_5, msg_to_check_it_18_cnu_52_in_0, msg_to_check_it_18_cnu_52_in_1, msg_to_check_it_18_cnu_52_in_2, msg_to_check_it_18_cnu_52_in_3, msg_to_check_it_18_cnu_52_in_4, msg_to_check_it_18_cnu_52_in_5, msg_to_check_it_18_cnu_53_in_0, msg_to_check_it_18_cnu_53_in_1, msg_to_check_it_18_cnu_53_in_2, msg_to_check_it_18_cnu_53_in_3, msg_to_check_it_18_cnu_53_in_4, msg_to_check_it_18_cnu_53_in_5, msg_to_check_it_18_cnu_54_in_0, msg_to_check_it_18_cnu_54_in_1, msg_to_check_it_18_cnu_54_in_2, msg_to_check_it_18_cnu_54_in_3, msg_to_check_it_18_cnu_54_in_4, msg_to_check_it_18_cnu_54_in_5, msg_to_check_it_18_cnu_55_in_0, msg_to_check_it_18_cnu_55_in_1, msg_to_check_it_18_cnu_55_in_2, msg_to_check_it_18_cnu_55_in_3, msg_to_check_it_18_cnu_55_in_4, msg_to_check_it_18_cnu_55_in_5, msg_to_check_it_18_cnu_56_in_0, msg_to_check_it_18_cnu_56_in_1, msg_to_check_it_18_cnu_56_in_2, msg_to_check_it_18_cnu_56_in_3, msg_to_check_it_18_cnu_56_in_4, msg_to_check_it_18_cnu_56_in_5, msg_to_check_it_18_cnu_57_in_0, msg_to_check_it_18_cnu_57_in_1, msg_to_check_it_18_cnu_57_in_2, msg_to_check_it_18_cnu_57_in_3, msg_to_check_it_18_cnu_57_in_4, msg_to_check_it_18_cnu_57_in_5, msg_to_check_it_18_cnu_58_in_0, msg_to_check_it_18_cnu_58_in_1, msg_to_check_it_18_cnu_58_in_2, msg_to_check_it_18_cnu_58_in_3, msg_to_check_it_18_cnu_58_in_4, msg_to_check_it_18_cnu_58_in_5, msg_to_check_it_18_cnu_59_in_0, msg_to_check_it_18_cnu_59_in_1, msg_to_check_it_18_cnu_59_in_2, msg_to_check_it_18_cnu_59_in_3, msg_to_check_it_18_cnu_59_in_4, msg_to_check_it_18_cnu_59_in_5, msg_to_check_it_18_cnu_60_in_0, msg_to_check_it_18_cnu_60_in_1, msg_to_check_it_18_cnu_60_in_2, msg_to_check_it_18_cnu_60_in_3, msg_to_check_it_18_cnu_60_in_4, msg_to_check_it_18_cnu_60_in_5, msg_to_check_it_18_cnu_61_in_0, msg_to_check_it_18_cnu_61_in_1, msg_to_check_it_18_cnu_61_in_2, msg_to_check_it_18_cnu_61_in_3, msg_to_check_it_18_cnu_61_in_4, msg_to_check_it_18_cnu_61_in_5, msg_to_check_it_18_cnu_62_in_0, msg_to_check_it_18_cnu_62_in_1, msg_to_check_it_18_cnu_62_in_2, msg_to_check_it_18_cnu_62_in_3, msg_to_check_it_18_cnu_62_in_4, msg_to_check_it_18_cnu_62_in_5, msg_to_check_it_18_cnu_63_in_0, msg_to_check_it_18_cnu_63_in_1, msg_to_check_it_18_cnu_63_in_2, msg_to_check_it_18_cnu_63_in_3, msg_to_check_it_18_cnu_63_in_4, msg_to_check_it_18_cnu_63_in_5, msg_to_check_it_18_cnu_64_in_0, msg_to_check_it_18_cnu_64_in_1, msg_to_check_it_18_cnu_64_in_2, msg_to_check_it_18_cnu_64_in_3, msg_to_check_it_18_cnu_64_in_4, msg_to_check_it_18_cnu_64_in_5, msg_to_check_it_18_cnu_65_in_0, msg_to_check_it_18_cnu_65_in_1, msg_to_check_it_18_cnu_65_in_2, msg_to_check_it_18_cnu_65_in_3, msg_to_check_it_18_cnu_65_in_4, msg_to_check_it_18_cnu_65_in_5, msg_to_check_it_18_cnu_66_in_0, msg_to_check_it_18_cnu_66_in_1, msg_to_check_it_18_cnu_66_in_2, msg_to_check_it_18_cnu_66_in_3, msg_to_check_it_18_cnu_66_in_4, msg_to_check_it_18_cnu_66_in_5, msg_to_check_it_18_cnu_67_in_0, msg_to_check_it_18_cnu_67_in_1, msg_to_check_it_18_cnu_67_in_2, msg_to_check_it_18_cnu_67_in_3, msg_to_check_it_18_cnu_67_in_4, msg_to_check_it_18_cnu_67_in_5, msg_to_check_it_18_cnu_68_in_0, msg_to_check_it_18_cnu_68_in_1, msg_to_check_it_18_cnu_68_in_2, msg_to_check_it_18_cnu_68_in_3, msg_to_check_it_18_cnu_68_in_4, msg_to_check_it_18_cnu_68_in_5, msg_to_check_it_18_cnu_69_in_0, msg_to_check_it_18_cnu_69_in_1, msg_to_check_it_18_cnu_69_in_2, msg_to_check_it_18_cnu_69_in_3, msg_to_check_it_18_cnu_69_in_4, msg_to_check_it_18_cnu_69_in_5, msg_to_check_it_18_cnu_70_in_0, msg_to_check_it_18_cnu_70_in_1, msg_to_check_it_18_cnu_70_in_2, msg_to_check_it_18_cnu_70_in_3, msg_to_check_it_18_cnu_70_in_4, msg_to_check_it_18_cnu_70_in_5, msg_to_check_it_18_cnu_71_in_0, msg_to_check_it_18_cnu_71_in_1, msg_to_check_it_18_cnu_71_in_2, msg_to_check_it_18_cnu_71_in_3, msg_to_check_it_18_cnu_71_in_4, msg_to_check_it_18_cnu_71_in_5, msg_to_check_it_18_cnu_72_in_0, msg_to_check_it_18_cnu_72_in_1, msg_to_check_it_18_cnu_72_in_2, msg_to_check_it_18_cnu_72_in_3, msg_to_check_it_18_cnu_72_in_4, msg_to_check_it_18_cnu_72_in_5, msg_to_check_it_18_cnu_73_in_0, msg_to_check_it_18_cnu_73_in_1, msg_to_check_it_18_cnu_73_in_2, msg_to_check_it_18_cnu_73_in_3, msg_to_check_it_18_cnu_73_in_4, msg_to_check_it_18_cnu_73_in_5, msg_to_check_it_18_cnu_74_in_0, msg_to_check_it_18_cnu_74_in_1, msg_to_check_it_18_cnu_74_in_2, msg_to_check_it_18_cnu_74_in_3, msg_to_check_it_18_cnu_74_in_4, msg_to_check_it_18_cnu_74_in_5, msg_to_check_it_18_cnu_75_in_0, msg_to_check_it_18_cnu_75_in_1, msg_to_check_it_18_cnu_75_in_2, msg_to_check_it_18_cnu_75_in_3, msg_to_check_it_18_cnu_75_in_4, msg_to_check_it_18_cnu_75_in_5, msg_to_check_it_18_cnu_76_in_0, msg_to_check_it_18_cnu_76_in_1, msg_to_check_it_18_cnu_76_in_2, msg_to_check_it_18_cnu_76_in_3, msg_to_check_it_18_cnu_76_in_4, msg_to_check_it_18_cnu_76_in_5, msg_to_check_it_18_cnu_77_in_0, msg_to_check_it_18_cnu_77_in_1, msg_to_check_it_18_cnu_77_in_2, msg_to_check_it_18_cnu_77_in_3, msg_to_check_it_18_cnu_77_in_4, msg_to_check_it_18_cnu_77_in_5, msg_to_check_it_18_cnu_78_in_0, msg_to_check_it_18_cnu_78_in_1, msg_to_check_it_18_cnu_78_in_2, msg_to_check_it_18_cnu_78_in_3, msg_to_check_it_18_cnu_78_in_4, msg_to_check_it_18_cnu_78_in_5, msg_to_check_it_18_cnu_79_in_0, msg_to_check_it_18_cnu_79_in_1, msg_to_check_it_18_cnu_79_in_2, msg_to_check_it_18_cnu_79_in_3, msg_to_check_it_18_cnu_79_in_4, msg_to_check_it_18_cnu_79_in_5, msg_to_check_it_18_cnu_80_in_0, msg_to_check_it_18_cnu_80_in_1, msg_to_check_it_18_cnu_80_in_2, msg_to_check_it_18_cnu_80_in_3, msg_to_check_it_18_cnu_80_in_4, msg_to_check_it_18_cnu_80_in_5, msg_to_check_it_18_cnu_81_in_0, msg_to_check_it_18_cnu_81_in_1, msg_to_check_it_18_cnu_81_in_2, msg_to_check_it_18_cnu_81_in_3, msg_to_check_it_18_cnu_81_in_4, msg_to_check_it_18_cnu_81_in_5, msg_to_check_it_18_cnu_82_in_0, msg_to_check_it_18_cnu_82_in_1, msg_to_check_it_18_cnu_82_in_2, msg_to_check_it_18_cnu_82_in_3, msg_to_check_it_18_cnu_82_in_4, msg_to_check_it_18_cnu_82_in_5, msg_to_check_it_18_cnu_83_in_0, msg_to_check_it_18_cnu_83_in_1, msg_to_check_it_18_cnu_83_in_2, msg_to_check_it_18_cnu_83_in_3, msg_to_check_it_18_cnu_83_in_4, msg_to_check_it_18_cnu_83_in_5, msg_to_check_it_18_cnu_84_in_0, msg_to_check_it_18_cnu_84_in_1, msg_to_check_it_18_cnu_84_in_2, msg_to_check_it_18_cnu_84_in_3, msg_to_check_it_18_cnu_84_in_4, msg_to_check_it_18_cnu_84_in_5, msg_to_check_it_18_cnu_85_in_0, msg_to_check_it_18_cnu_85_in_1, msg_to_check_it_18_cnu_85_in_2, msg_to_check_it_18_cnu_85_in_3, msg_to_check_it_18_cnu_85_in_4, msg_to_check_it_18_cnu_85_in_5, msg_to_check_it_18_cnu_86_in_0, msg_to_check_it_18_cnu_86_in_1, msg_to_check_it_18_cnu_86_in_2, msg_to_check_it_18_cnu_86_in_3, msg_to_check_it_18_cnu_86_in_4, msg_to_check_it_18_cnu_86_in_5, msg_to_check_it_18_cnu_87_in_0, msg_to_check_it_18_cnu_87_in_1, msg_to_check_it_18_cnu_87_in_2, msg_to_check_it_18_cnu_87_in_3, msg_to_check_it_18_cnu_87_in_4, msg_to_check_it_18_cnu_87_in_5, msg_to_check_it_18_cnu_88_in_0, msg_to_check_it_18_cnu_88_in_1, msg_to_check_it_18_cnu_88_in_2, msg_to_check_it_18_cnu_88_in_3, msg_to_check_it_18_cnu_88_in_4, msg_to_check_it_18_cnu_88_in_5, msg_to_check_it_18_cnu_89_in_0, msg_to_check_it_18_cnu_89_in_1, msg_to_check_it_18_cnu_89_in_2, msg_to_check_it_18_cnu_89_in_3, msg_to_check_it_18_cnu_89_in_4, msg_to_check_it_18_cnu_89_in_5, msg_to_check_it_18_cnu_90_in_0, msg_to_check_it_18_cnu_90_in_1, msg_to_check_it_18_cnu_90_in_2, msg_to_check_it_18_cnu_90_in_3, msg_to_check_it_18_cnu_90_in_4, msg_to_check_it_18_cnu_90_in_5, msg_to_check_it_18_cnu_91_in_0, msg_to_check_it_18_cnu_91_in_1, msg_to_check_it_18_cnu_91_in_2, msg_to_check_it_18_cnu_91_in_3, msg_to_check_it_18_cnu_91_in_4, msg_to_check_it_18_cnu_91_in_5, msg_to_check_it_18_cnu_92_in_0, msg_to_check_it_18_cnu_92_in_1, msg_to_check_it_18_cnu_92_in_2, msg_to_check_it_18_cnu_92_in_3, msg_to_check_it_18_cnu_92_in_4, msg_to_check_it_18_cnu_92_in_5, msg_to_check_it_18_cnu_93_in_0, msg_to_check_it_18_cnu_93_in_1, msg_to_check_it_18_cnu_93_in_2, msg_to_check_it_18_cnu_93_in_3, msg_to_check_it_18_cnu_93_in_4, msg_to_check_it_18_cnu_93_in_5, msg_to_check_it_18_cnu_94_in_0, msg_to_check_it_18_cnu_94_in_1, msg_to_check_it_18_cnu_94_in_2, msg_to_check_it_18_cnu_94_in_3, msg_to_check_it_18_cnu_94_in_4, msg_to_check_it_18_cnu_94_in_5, msg_to_check_it_18_cnu_95_in_0, msg_to_check_it_18_cnu_95_in_1, msg_to_check_it_18_cnu_95_in_2, msg_to_check_it_18_cnu_95_in_3, msg_to_check_it_18_cnu_95_in_4, msg_to_check_it_18_cnu_95_in_5, msg_to_check_it_18_cnu_96_in_0, msg_to_check_it_18_cnu_96_in_1, msg_to_check_it_18_cnu_96_in_2, msg_to_check_it_18_cnu_96_in_3, msg_to_check_it_18_cnu_96_in_4, msg_to_check_it_18_cnu_96_in_5, msg_to_check_it_18_cnu_97_in_0, msg_to_check_it_18_cnu_97_in_1, msg_to_check_it_18_cnu_97_in_2, msg_to_check_it_18_cnu_97_in_3, msg_to_check_it_18_cnu_97_in_4, msg_to_check_it_18_cnu_97_in_5, msg_to_check_it_18_cnu_98_in_0, msg_to_check_it_18_cnu_98_in_1, msg_to_check_it_18_cnu_98_in_2, msg_to_check_it_18_cnu_98_in_3, msg_to_check_it_18_cnu_98_in_4, msg_to_check_it_18_cnu_98_in_5, msg_to_check_it_19_cnu_0_in_0, msg_to_check_it_19_cnu_0_in_1, msg_to_check_it_19_cnu_0_in_2, msg_to_check_it_19_cnu_0_in_3, msg_to_check_it_19_cnu_0_in_4, msg_to_check_it_19_cnu_0_in_5, msg_to_check_it_19_cnu_1_in_0, msg_to_check_it_19_cnu_1_in_1, msg_to_check_it_19_cnu_1_in_2, msg_to_check_it_19_cnu_1_in_3, msg_to_check_it_19_cnu_1_in_4, msg_to_check_it_19_cnu_1_in_5, msg_to_check_it_19_cnu_2_in_0, msg_to_check_it_19_cnu_2_in_1, msg_to_check_it_19_cnu_2_in_2, msg_to_check_it_19_cnu_2_in_3, msg_to_check_it_19_cnu_2_in_4, msg_to_check_it_19_cnu_2_in_5, msg_to_check_it_19_cnu_3_in_0, msg_to_check_it_19_cnu_3_in_1, msg_to_check_it_19_cnu_3_in_2, msg_to_check_it_19_cnu_3_in_3, msg_to_check_it_19_cnu_3_in_4, msg_to_check_it_19_cnu_3_in_5, msg_to_check_it_19_cnu_4_in_0, msg_to_check_it_19_cnu_4_in_1, msg_to_check_it_19_cnu_4_in_2, msg_to_check_it_19_cnu_4_in_3, msg_to_check_it_19_cnu_4_in_4, msg_to_check_it_19_cnu_4_in_5, msg_to_check_it_19_cnu_5_in_0, msg_to_check_it_19_cnu_5_in_1, msg_to_check_it_19_cnu_5_in_2, msg_to_check_it_19_cnu_5_in_3, msg_to_check_it_19_cnu_5_in_4, msg_to_check_it_19_cnu_5_in_5, msg_to_check_it_19_cnu_6_in_0, msg_to_check_it_19_cnu_6_in_1, msg_to_check_it_19_cnu_6_in_2, msg_to_check_it_19_cnu_6_in_3, msg_to_check_it_19_cnu_6_in_4, msg_to_check_it_19_cnu_6_in_5, msg_to_check_it_19_cnu_7_in_0, msg_to_check_it_19_cnu_7_in_1, msg_to_check_it_19_cnu_7_in_2, msg_to_check_it_19_cnu_7_in_3, msg_to_check_it_19_cnu_7_in_4, msg_to_check_it_19_cnu_7_in_5, msg_to_check_it_19_cnu_8_in_0, msg_to_check_it_19_cnu_8_in_1, msg_to_check_it_19_cnu_8_in_2, msg_to_check_it_19_cnu_8_in_3, msg_to_check_it_19_cnu_8_in_4, msg_to_check_it_19_cnu_8_in_5, msg_to_check_it_19_cnu_9_in_0, msg_to_check_it_19_cnu_9_in_1, msg_to_check_it_19_cnu_9_in_2, msg_to_check_it_19_cnu_9_in_3, msg_to_check_it_19_cnu_9_in_4, msg_to_check_it_19_cnu_9_in_5, msg_to_check_it_19_cnu_10_in_0, msg_to_check_it_19_cnu_10_in_1, msg_to_check_it_19_cnu_10_in_2, msg_to_check_it_19_cnu_10_in_3, msg_to_check_it_19_cnu_10_in_4, msg_to_check_it_19_cnu_10_in_5, msg_to_check_it_19_cnu_11_in_0, msg_to_check_it_19_cnu_11_in_1, msg_to_check_it_19_cnu_11_in_2, msg_to_check_it_19_cnu_11_in_3, msg_to_check_it_19_cnu_11_in_4, msg_to_check_it_19_cnu_11_in_5, msg_to_check_it_19_cnu_12_in_0, msg_to_check_it_19_cnu_12_in_1, msg_to_check_it_19_cnu_12_in_2, msg_to_check_it_19_cnu_12_in_3, msg_to_check_it_19_cnu_12_in_4, msg_to_check_it_19_cnu_12_in_5, msg_to_check_it_19_cnu_13_in_0, msg_to_check_it_19_cnu_13_in_1, msg_to_check_it_19_cnu_13_in_2, msg_to_check_it_19_cnu_13_in_3, msg_to_check_it_19_cnu_13_in_4, msg_to_check_it_19_cnu_13_in_5, msg_to_check_it_19_cnu_14_in_0, msg_to_check_it_19_cnu_14_in_1, msg_to_check_it_19_cnu_14_in_2, msg_to_check_it_19_cnu_14_in_3, msg_to_check_it_19_cnu_14_in_4, msg_to_check_it_19_cnu_14_in_5, msg_to_check_it_19_cnu_15_in_0, msg_to_check_it_19_cnu_15_in_1, msg_to_check_it_19_cnu_15_in_2, msg_to_check_it_19_cnu_15_in_3, msg_to_check_it_19_cnu_15_in_4, msg_to_check_it_19_cnu_15_in_5, msg_to_check_it_19_cnu_16_in_0, msg_to_check_it_19_cnu_16_in_1, msg_to_check_it_19_cnu_16_in_2, msg_to_check_it_19_cnu_16_in_3, msg_to_check_it_19_cnu_16_in_4, msg_to_check_it_19_cnu_16_in_5, msg_to_check_it_19_cnu_17_in_0, msg_to_check_it_19_cnu_17_in_1, msg_to_check_it_19_cnu_17_in_2, msg_to_check_it_19_cnu_17_in_3, msg_to_check_it_19_cnu_17_in_4, msg_to_check_it_19_cnu_17_in_5, msg_to_check_it_19_cnu_18_in_0, msg_to_check_it_19_cnu_18_in_1, msg_to_check_it_19_cnu_18_in_2, msg_to_check_it_19_cnu_18_in_3, msg_to_check_it_19_cnu_18_in_4, msg_to_check_it_19_cnu_18_in_5, msg_to_check_it_19_cnu_19_in_0, msg_to_check_it_19_cnu_19_in_1, msg_to_check_it_19_cnu_19_in_2, msg_to_check_it_19_cnu_19_in_3, msg_to_check_it_19_cnu_19_in_4, msg_to_check_it_19_cnu_19_in_5, msg_to_check_it_19_cnu_20_in_0, msg_to_check_it_19_cnu_20_in_1, msg_to_check_it_19_cnu_20_in_2, msg_to_check_it_19_cnu_20_in_3, msg_to_check_it_19_cnu_20_in_4, msg_to_check_it_19_cnu_20_in_5, msg_to_check_it_19_cnu_21_in_0, msg_to_check_it_19_cnu_21_in_1, msg_to_check_it_19_cnu_21_in_2, msg_to_check_it_19_cnu_21_in_3, msg_to_check_it_19_cnu_21_in_4, msg_to_check_it_19_cnu_21_in_5, msg_to_check_it_19_cnu_22_in_0, msg_to_check_it_19_cnu_22_in_1, msg_to_check_it_19_cnu_22_in_2, msg_to_check_it_19_cnu_22_in_3, msg_to_check_it_19_cnu_22_in_4, msg_to_check_it_19_cnu_22_in_5, msg_to_check_it_19_cnu_23_in_0, msg_to_check_it_19_cnu_23_in_1, msg_to_check_it_19_cnu_23_in_2, msg_to_check_it_19_cnu_23_in_3, msg_to_check_it_19_cnu_23_in_4, msg_to_check_it_19_cnu_23_in_5, msg_to_check_it_19_cnu_24_in_0, msg_to_check_it_19_cnu_24_in_1, msg_to_check_it_19_cnu_24_in_2, msg_to_check_it_19_cnu_24_in_3, msg_to_check_it_19_cnu_24_in_4, msg_to_check_it_19_cnu_24_in_5, msg_to_check_it_19_cnu_25_in_0, msg_to_check_it_19_cnu_25_in_1, msg_to_check_it_19_cnu_25_in_2, msg_to_check_it_19_cnu_25_in_3, msg_to_check_it_19_cnu_25_in_4, msg_to_check_it_19_cnu_25_in_5, msg_to_check_it_19_cnu_26_in_0, msg_to_check_it_19_cnu_26_in_1, msg_to_check_it_19_cnu_26_in_2, msg_to_check_it_19_cnu_26_in_3, msg_to_check_it_19_cnu_26_in_4, msg_to_check_it_19_cnu_26_in_5, msg_to_check_it_19_cnu_27_in_0, msg_to_check_it_19_cnu_27_in_1, msg_to_check_it_19_cnu_27_in_2, msg_to_check_it_19_cnu_27_in_3, msg_to_check_it_19_cnu_27_in_4, msg_to_check_it_19_cnu_27_in_5, msg_to_check_it_19_cnu_28_in_0, msg_to_check_it_19_cnu_28_in_1, msg_to_check_it_19_cnu_28_in_2, msg_to_check_it_19_cnu_28_in_3, msg_to_check_it_19_cnu_28_in_4, msg_to_check_it_19_cnu_28_in_5, msg_to_check_it_19_cnu_29_in_0, msg_to_check_it_19_cnu_29_in_1, msg_to_check_it_19_cnu_29_in_2, msg_to_check_it_19_cnu_29_in_3, msg_to_check_it_19_cnu_29_in_4, msg_to_check_it_19_cnu_29_in_5, msg_to_check_it_19_cnu_30_in_0, msg_to_check_it_19_cnu_30_in_1, msg_to_check_it_19_cnu_30_in_2, msg_to_check_it_19_cnu_30_in_3, msg_to_check_it_19_cnu_30_in_4, msg_to_check_it_19_cnu_30_in_5, msg_to_check_it_19_cnu_31_in_0, msg_to_check_it_19_cnu_31_in_1, msg_to_check_it_19_cnu_31_in_2, msg_to_check_it_19_cnu_31_in_3, msg_to_check_it_19_cnu_31_in_4, msg_to_check_it_19_cnu_31_in_5, msg_to_check_it_19_cnu_32_in_0, msg_to_check_it_19_cnu_32_in_1, msg_to_check_it_19_cnu_32_in_2, msg_to_check_it_19_cnu_32_in_3, msg_to_check_it_19_cnu_32_in_4, msg_to_check_it_19_cnu_32_in_5, msg_to_check_it_19_cnu_33_in_0, msg_to_check_it_19_cnu_33_in_1, msg_to_check_it_19_cnu_33_in_2, msg_to_check_it_19_cnu_33_in_3, msg_to_check_it_19_cnu_33_in_4, msg_to_check_it_19_cnu_33_in_5, msg_to_check_it_19_cnu_34_in_0, msg_to_check_it_19_cnu_34_in_1, msg_to_check_it_19_cnu_34_in_2, msg_to_check_it_19_cnu_34_in_3, msg_to_check_it_19_cnu_34_in_4, msg_to_check_it_19_cnu_34_in_5, msg_to_check_it_19_cnu_35_in_0, msg_to_check_it_19_cnu_35_in_1, msg_to_check_it_19_cnu_35_in_2, msg_to_check_it_19_cnu_35_in_3, msg_to_check_it_19_cnu_35_in_4, msg_to_check_it_19_cnu_35_in_5, msg_to_check_it_19_cnu_36_in_0, msg_to_check_it_19_cnu_36_in_1, msg_to_check_it_19_cnu_36_in_2, msg_to_check_it_19_cnu_36_in_3, msg_to_check_it_19_cnu_36_in_4, msg_to_check_it_19_cnu_36_in_5, msg_to_check_it_19_cnu_37_in_0, msg_to_check_it_19_cnu_37_in_1, msg_to_check_it_19_cnu_37_in_2, msg_to_check_it_19_cnu_37_in_3, msg_to_check_it_19_cnu_37_in_4, msg_to_check_it_19_cnu_37_in_5, msg_to_check_it_19_cnu_38_in_0, msg_to_check_it_19_cnu_38_in_1, msg_to_check_it_19_cnu_38_in_2, msg_to_check_it_19_cnu_38_in_3, msg_to_check_it_19_cnu_38_in_4, msg_to_check_it_19_cnu_38_in_5, msg_to_check_it_19_cnu_39_in_0, msg_to_check_it_19_cnu_39_in_1, msg_to_check_it_19_cnu_39_in_2, msg_to_check_it_19_cnu_39_in_3, msg_to_check_it_19_cnu_39_in_4, msg_to_check_it_19_cnu_39_in_5, msg_to_check_it_19_cnu_40_in_0, msg_to_check_it_19_cnu_40_in_1, msg_to_check_it_19_cnu_40_in_2, msg_to_check_it_19_cnu_40_in_3, msg_to_check_it_19_cnu_40_in_4, msg_to_check_it_19_cnu_40_in_5, msg_to_check_it_19_cnu_41_in_0, msg_to_check_it_19_cnu_41_in_1, msg_to_check_it_19_cnu_41_in_2, msg_to_check_it_19_cnu_41_in_3, msg_to_check_it_19_cnu_41_in_4, msg_to_check_it_19_cnu_41_in_5, msg_to_check_it_19_cnu_42_in_0, msg_to_check_it_19_cnu_42_in_1, msg_to_check_it_19_cnu_42_in_2, msg_to_check_it_19_cnu_42_in_3, msg_to_check_it_19_cnu_42_in_4, msg_to_check_it_19_cnu_42_in_5, msg_to_check_it_19_cnu_43_in_0, msg_to_check_it_19_cnu_43_in_1, msg_to_check_it_19_cnu_43_in_2, msg_to_check_it_19_cnu_43_in_3, msg_to_check_it_19_cnu_43_in_4, msg_to_check_it_19_cnu_43_in_5, msg_to_check_it_19_cnu_44_in_0, msg_to_check_it_19_cnu_44_in_1, msg_to_check_it_19_cnu_44_in_2, msg_to_check_it_19_cnu_44_in_3, msg_to_check_it_19_cnu_44_in_4, msg_to_check_it_19_cnu_44_in_5, msg_to_check_it_19_cnu_45_in_0, msg_to_check_it_19_cnu_45_in_1, msg_to_check_it_19_cnu_45_in_2, msg_to_check_it_19_cnu_45_in_3, msg_to_check_it_19_cnu_45_in_4, msg_to_check_it_19_cnu_45_in_5, msg_to_check_it_19_cnu_46_in_0, msg_to_check_it_19_cnu_46_in_1, msg_to_check_it_19_cnu_46_in_2, msg_to_check_it_19_cnu_46_in_3, msg_to_check_it_19_cnu_46_in_4, msg_to_check_it_19_cnu_46_in_5, msg_to_check_it_19_cnu_47_in_0, msg_to_check_it_19_cnu_47_in_1, msg_to_check_it_19_cnu_47_in_2, msg_to_check_it_19_cnu_47_in_3, msg_to_check_it_19_cnu_47_in_4, msg_to_check_it_19_cnu_47_in_5, msg_to_check_it_19_cnu_48_in_0, msg_to_check_it_19_cnu_48_in_1, msg_to_check_it_19_cnu_48_in_2, msg_to_check_it_19_cnu_48_in_3, msg_to_check_it_19_cnu_48_in_4, msg_to_check_it_19_cnu_48_in_5, msg_to_check_it_19_cnu_49_in_0, msg_to_check_it_19_cnu_49_in_1, msg_to_check_it_19_cnu_49_in_2, msg_to_check_it_19_cnu_49_in_3, msg_to_check_it_19_cnu_49_in_4, msg_to_check_it_19_cnu_49_in_5, msg_to_check_it_19_cnu_50_in_0, msg_to_check_it_19_cnu_50_in_1, msg_to_check_it_19_cnu_50_in_2, msg_to_check_it_19_cnu_50_in_3, msg_to_check_it_19_cnu_50_in_4, msg_to_check_it_19_cnu_50_in_5, msg_to_check_it_19_cnu_51_in_0, msg_to_check_it_19_cnu_51_in_1, msg_to_check_it_19_cnu_51_in_2, msg_to_check_it_19_cnu_51_in_3, msg_to_check_it_19_cnu_51_in_4, msg_to_check_it_19_cnu_51_in_5, msg_to_check_it_19_cnu_52_in_0, msg_to_check_it_19_cnu_52_in_1, msg_to_check_it_19_cnu_52_in_2, msg_to_check_it_19_cnu_52_in_3, msg_to_check_it_19_cnu_52_in_4, msg_to_check_it_19_cnu_52_in_5, msg_to_check_it_19_cnu_53_in_0, msg_to_check_it_19_cnu_53_in_1, msg_to_check_it_19_cnu_53_in_2, msg_to_check_it_19_cnu_53_in_3, msg_to_check_it_19_cnu_53_in_4, msg_to_check_it_19_cnu_53_in_5, msg_to_check_it_19_cnu_54_in_0, msg_to_check_it_19_cnu_54_in_1, msg_to_check_it_19_cnu_54_in_2, msg_to_check_it_19_cnu_54_in_3, msg_to_check_it_19_cnu_54_in_4, msg_to_check_it_19_cnu_54_in_5, msg_to_check_it_19_cnu_55_in_0, msg_to_check_it_19_cnu_55_in_1, msg_to_check_it_19_cnu_55_in_2, msg_to_check_it_19_cnu_55_in_3, msg_to_check_it_19_cnu_55_in_4, msg_to_check_it_19_cnu_55_in_5, msg_to_check_it_19_cnu_56_in_0, msg_to_check_it_19_cnu_56_in_1, msg_to_check_it_19_cnu_56_in_2, msg_to_check_it_19_cnu_56_in_3, msg_to_check_it_19_cnu_56_in_4, msg_to_check_it_19_cnu_56_in_5, msg_to_check_it_19_cnu_57_in_0, msg_to_check_it_19_cnu_57_in_1, msg_to_check_it_19_cnu_57_in_2, msg_to_check_it_19_cnu_57_in_3, msg_to_check_it_19_cnu_57_in_4, msg_to_check_it_19_cnu_57_in_5, msg_to_check_it_19_cnu_58_in_0, msg_to_check_it_19_cnu_58_in_1, msg_to_check_it_19_cnu_58_in_2, msg_to_check_it_19_cnu_58_in_3, msg_to_check_it_19_cnu_58_in_4, msg_to_check_it_19_cnu_58_in_5, msg_to_check_it_19_cnu_59_in_0, msg_to_check_it_19_cnu_59_in_1, msg_to_check_it_19_cnu_59_in_2, msg_to_check_it_19_cnu_59_in_3, msg_to_check_it_19_cnu_59_in_4, msg_to_check_it_19_cnu_59_in_5, msg_to_check_it_19_cnu_60_in_0, msg_to_check_it_19_cnu_60_in_1, msg_to_check_it_19_cnu_60_in_2, msg_to_check_it_19_cnu_60_in_3, msg_to_check_it_19_cnu_60_in_4, msg_to_check_it_19_cnu_60_in_5, msg_to_check_it_19_cnu_61_in_0, msg_to_check_it_19_cnu_61_in_1, msg_to_check_it_19_cnu_61_in_2, msg_to_check_it_19_cnu_61_in_3, msg_to_check_it_19_cnu_61_in_4, msg_to_check_it_19_cnu_61_in_5, msg_to_check_it_19_cnu_62_in_0, msg_to_check_it_19_cnu_62_in_1, msg_to_check_it_19_cnu_62_in_2, msg_to_check_it_19_cnu_62_in_3, msg_to_check_it_19_cnu_62_in_4, msg_to_check_it_19_cnu_62_in_5, msg_to_check_it_19_cnu_63_in_0, msg_to_check_it_19_cnu_63_in_1, msg_to_check_it_19_cnu_63_in_2, msg_to_check_it_19_cnu_63_in_3, msg_to_check_it_19_cnu_63_in_4, msg_to_check_it_19_cnu_63_in_5, msg_to_check_it_19_cnu_64_in_0, msg_to_check_it_19_cnu_64_in_1, msg_to_check_it_19_cnu_64_in_2, msg_to_check_it_19_cnu_64_in_3, msg_to_check_it_19_cnu_64_in_4, msg_to_check_it_19_cnu_64_in_5, msg_to_check_it_19_cnu_65_in_0, msg_to_check_it_19_cnu_65_in_1, msg_to_check_it_19_cnu_65_in_2, msg_to_check_it_19_cnu_65_in_3, msg_to_check_it_19_cnu_65_in_4, msg_to_check_it_19_cnu_65_in_5, msg_to_check_it_19_cnu_66_in_0, msg_to_check_it_19_cnu_66_in_1, msg_to_check_it_19_cnu_66_in_2, msg_to_check_it_19_cnu_66_in_3, msg_to_check_it_19_cnu_66_in_4, msg_to_check_it_19_cnu_66_in_5, msg_to_check_it_19_cnu_67_in_0, msg_to_check_it_19_cnu_67_in_1, msg_to_check_it_19_cnu_67_in_2, msg_to_check_it_19_cnu_67_in_3, msg_to_check_it_19_cnu_67_in_4, msg_to_check_it_19_cnu_67_in_5, msg_to_check_it_19_cnu_68_in_0, msg_to_check_it_19_cnu_68_in_1, msg_to_check_it_19_cnu_68_in_2, msg_to_check_it_19_cnu_68_in_3, msg_to_check_it_19_cnu_68_in_4, msg_to_check_it_19_cnu_68_in_5, msg_to_check_it_19_cnu_69_in_0, msg_to_check_it_19_cnu_69_in_1, msg_to_check_it_19_cnu_69_in_2, msg_to_check_it_19_cnu_69_in_3, msg_to_check_it_19_cnu_69_in_4, msg_to_check_it_19_cnu_69_in_5, msg_to_check_it_19_cnu_70_in_0, msg_to_check_it_19_cnu_70_in_1, msg_to_check_it_19_cnu_70_in_2, msg_to_check_it_19_cnu_70_in_3, msg_to_check_it_19_cnu_70_in_4, msg_to_check_it_19_cnu_70_in_5, msg_to_check_it_19_cnu_71_in_0, msg_to_check_it_19_cnu_71_in_1, msg_to_check_it_19_cnu_71_in_2, msg_to_check_it_19_cnu_71_in_3, msg_to_check_it_19_cnu_71_in_4, msg_to_check_it_19_cnu_71_in_5, msg_to_check_it_19_cnu_72_in_0, msg_to_check_it_19_cnu_72_in_1, msg_to_check_it_19_cnu_72_in_2, msg_to_check_it_19_cnu_72_in_3, msg_to_check_it_19_cnu_72_in_4, msg_to_check_it_19_cnu_72_in_5, msg_to_check_it_19_cnu_73_in_0, msg_to_check_it_19_cnu_73_in_1, msg_to_check_it_19_cnu_73_in_2, msg_to_check_it_19_cnu_73_in_3, msg_to_check_it_19_cnu_73_in_4, msg_to_check_it_19_cnu_73_in_5, msg_to_check_it_19_cnu_74_in_0, msg_to_check_it_19_cnu_74_in_1, msg_to_check_it_19_cnu_74_in_2, msg_to_check_it_19_cnu_74_in_3, msg_to_check_it_19_cnu_74_in_4, msg_to_check_it_19_cnu_74_in_5, msg_to_check_it_19_cnu_75_in_0, msg_to_check_it_19_cnu_75_in_1, msg_to_check_it_19_cnu_75_in_2, msg_to_check_it_19_cnu_75_in_3, msg_to_check_it_19_cnu_75_in_4, msg_to_check_it_19_cnu_75_in_5, msg_to_check_it_19_cnu_76_in_0, msg_to_check_it_19_cnu_76_in_1, msg_to_check_it_19_cnu_76_in_2, msg_to_check_it_19_cnu_76_in_3, msg_to_check_it_19_cnu_76_in_4, msg_to_check_it_19_cnu_76_in_5, msg_to_check_it_19_cnu_77_in_0, msg_to_check_it_19_cnu_77_in_1, msg_to_check_it_19_cnu_77_in_2, msg_to_check_it_19_cnu_77_in_3, msg_to_check_it_19_cnu_77_in_4, msg_to_check_it_19_cnu_77_in_5, msg_to_check_it_19_cnu_78_in_0, msg_to_check_it_19_cnu_78_in_1, msg_to_check_it_19_cnu_78_in_2, msg_to_check_it_19_cnu_78_in_3, msg_to_check_it_19_cnu_78_in_4, msg_to_check_it_19_cnu_78_in_5, msg_to_check_it_19_cnu_79_in_0, msg_to_check_it_19_cnu_79_in_1, msg_to_check_it_19_cnu_79_in_2, msg_to_check_it_19_cnu_79_in_3, msg_to_check_it_19_cnu_79_in_4, msg_to_check_it_19_cnu_79_in_5, msg_to_check_it_19_cnu_80_in_0, msg_to_check_it_19_cnu_80_in_1, msg_to_check_it_19_cnu_80_in_2, msg_to_check_it_19_cnu_80_in_3, msg_to_check_it_19_cnu_80_in_4, msg_to_check_it_19_cnu_80_in_5, msg_to_check_it_19_cnu_81_in_0, msg_to_check_it_19_cnu_81_in_1, msg_to_check_it_19_cnu_81_in_2, msg_to_check_it_19_cnu_81_in_3, msg_to_check_it_19_cnu_81_in_4, msg_to_check_it_19_cnu_81_in_5, msg_to_check_it_19_cnu_82_in_0, msg_to_check_it_19_cnu_82_in_1, msg_to_check_it_19_cnu_82_in_2, msg_to_check_it_19_cnu_82_in_3, msg_to_check_it_19_cnu_82_in_4, msg_to_check_it_19_cnu_82_in_5, msg_to_check_it_19_cnu_83_in_0, msg_to_check_it_19_cnu_83_in_1, msg_to_check_it_19_cnu_83_in_2, msg_to_check_it_19_cnu_83_in_3, msg_to_check_it_19_cnu_83_in_4, msg_to_check_it_19_cnu_83_in_5, msg_to_check_it_19_cnu_84_in_0, msg_to_check_it_19_cnu_84_in_1, msg_to_check_it_19_cnu_84_in_2, msg_to_check_it_19_cnu_84_in_3, msg_to_check_it_19_cnu_84_in_4, msg_to_check_it_19_cnu_84_in_5, msg_to_check_it_19_cnu_85_in_0, msg_to_check_it_19_cnu_85_in_1, msg_to_check_it_19_cnu_85_in_2, msg_to_check_it_19_cnu_85_in_3, msg_to_check_it_19_cnu_85_in_4, msg_to_check_it_19_cnu_85_in_5, msg_to_check_it_19_cnu_86_in_0, msg_to_check_it_19_cnu_86_in_1, msg_to_check_it_19_cnu_86_in_2, msg_to_check_it_19_cnu_86_in_3, msg_to_check_it_19_cnu_86_in_4, msg_to_check_it_19_cnu_86_in_5, msg_to_check_it_19_cnu_87_in_0, msg_to_check_it_19_cnu_87_in_1, msg_to_check_it_19_cnu_87_in_2, msg_to_check_it_19_cnu_87_in_3, msg_to_check_it_19_cnu_87_in_4, msg_to_check_it_19_cnu_87_in_5, msg_to_check_it_19_cnu_88_in_0, msg_to_check_it_19_cnu_88_in_1, msg_to_check_it_19_cnu_88_in_2, msg_to_check_it_19_cnu_88_in_3, msg_to_check_it_19_cnu_88_in_4, msg_to_check_it_19_cnu_88_in_5, msg_to_check_it_19_cnu_89_in_0, msg_to_check_it_19_cnu_89_in_1, msg_to_check_it_19_cnu_89_in_2, msg_to_check_it_19_cnu_89_in_3, msg_to_check_it_19_cnu_89_in_4, msg_to_check_it_19_cnu_89_in_5, msg_to_check_it_19_cnu_90_in_0, msg_to_check_it_19_cnu_90_in_1, msg_to_check_it_19_cnu_90_in_2, msg_to_check_it_19_cnu_90_in_3, msg_to_check_it_19_cnu_90_in_4, msg_to_check_it_19_cnu_90_in_5, msg_to_check_it_19_cnu_91_in_0, msg_to_check_it_19_cnu_91_in_1, msg_to_check_it_19_cnu_91_in_2, msg_to_check_it_19_cnu_91_in_3, msg_to_check_it_19_cnu_91_in_4, msg_to_check_it_19_cnu_91_in_5, msg_to_check_it_19_cnu_92_in_0, msg_to_check_it_19_cnu_92_in_1, msg_to_check_it_19_cnu_92_in_2, msg_to_check_it_19_cnu_92_in_3, msg_to_check_it_19_cnu_92_in_4, msg_to_check_it_19_cnu_92_in_5, msg_to_check_it_19_cnu_93_in_0, msg_to_check_it_19_cnu_93_in_1, msg_to_check_it_19_cnu_93_in_2, msg_to_check_it_19_cnu_93_in_3, msg_to_check_it_19_cnu_93_in_4, msg_to_check_it_19_cnu_93_in_5, msg_to_check_it_19_cnu_94_in_0, msg_to_check_it_19_cnu_94_in_1, msg_to_check_it_19_cnu_94_in_2, msg_to_check_it_19_cnu_94_in_3, msg_to_check_it_19_cnu_94_in_4, msg_to_check_it_19_cnu_94_in_5, msg_to_check_it_19_cnu_95_in_0, msg_to_check_it_19_cnu_95_in_1, msg_to_check_it_19_cnu_95_in_2, msg_to_check_it_19_cnu_95_in_3, msg_to_check_it_19_cnu_95_in_4, msg_to_check_it_19_cnu_95_in_5, msg_to_check_it_19_cnu_96_in_0, msg_to_check_it_19_cnu_96_in_1, msg_to_check_it_19_cnu_96_in_2, msg_to_check_it_19_cnu_96_in_3, msg_to_check_it_19_cnu_96_in_4, msg_to_check_it_19_cnu_96_in_5, msg_to_check_it_19_cnu_97_in_0, msg_to_check_it_19_cnu_97_in_1, msg_to_check_it_19_cnu_97_in_2, msg_to_check_it_19_cnu_97_in_3, msg_to_check_it_19_cnu_97_in_4, msg_to_check_it_19_cnu_97_in_5, msg_to_check_it_19_cnu_98_in_0, msg_to_check_it_19_cnu_98_in_1, msg_to_check_it_19_cnu_98_in_2, msg_to_check_it_19_cnu_98_in_3, msg_to_check_it_19_cnu_98_in_4, msg_to_check_it_19_cnu_98_in_5;
wire [7:0] msg_to_bit_it_1_vnu_0_in_0, msg_to_bit_it_1_vnu_0_in_1, msg_to_bit_it_1_vnu_0_in_2, msg_to_bit_it_1_vnu_1_in_0, msg_to_bit_it_1_vnu_1_in_1, msg_to_bit_it_1_vnu_1_in_2, msg_to_bit_it_1_vnu_2_in_0, msg_to_bit_it_1_vnu_2_in_1, msg_to_bit_it_1_vnu_2_in_2, msg_to_bit_it_1_vnu_3_in_0, msg_to_bit_it_1_vnu_3_in_1, msg_to_bit_it_1_vnu_3_in_2, msg_to_bit_it_1_vnu_4_in_0, msg_to_bit_it_1_vnu_4_in_1, msg_to_bit_it_1_vnu_4_in_2, msg_to_bit_it_1_vnu_5_in_0, msg_to_bit_it_1_vnu_5_in_1, msg_to_bit_it_1_vnu_5_in_2, msg_to_bit_it_1_vnu_6_in_0, msg_to_bit_it_1_vnu_6_in_1, msg_to_bit_it_1_vnu_6_in_2, msg_to_bit_it_1_vnu_7_in_0, msg_to_bit_it_1_vnu_7_in_1, msg_to_bit_it_1_vnu_7_in_2, msg_to_bit_it_1_vnu_8_in_0, msg_to_bit_it_1_vnu_8_in_1, msg_to_bit_it_1_vnu_8_in_2, msg_to_bit_it_1_vnu_9_in_0, msg_to_bit_it_1_vnu_9_in_1, msg_to_bit_it_1_vnu_9_in_2, msg_to_bit_it_1_vnu_10_in_0, msg_to_bit_it_1_vnu_10_in_1, msg_to_bit_it_1_vnu_10_in_2, msg_to_bit_it_1_vnu_11_in_0, msg_to_bit_it_1_vnu_11_in_1, msg_to_bit_it_1_vnu_11_in_2, msg_to_bit_it_1_vnu_12_in_0, msg_to_bit_it_1_vnu_12_in_1, msg_to_bit_it_1_vnu_12_in_2, msg_to_bit_it_1_vnu_13_in_0, msg_to_bit_it_1_vnu_13_in_1, msg_to_bit_it_1_vnu_13_in_2, msg_to_bit_it_1_vnu_14_in_0, msg_to_bit_it_1_vnu_14_in_1, msg_to_bit_it_1_vnu_14_in_2, msg_to_bit_it_1_vnu_15_in_0, msg_to_bit_it_1_vnu_15_in_1, msg_to_bit_it_1_vnu_15_in_2, msg_to_bit_it_1_vnu_16_in_0, msg_to_bit_it_1_vnu_16_in_1, msg_to_bit_it_1_vnu_16_in_2, msg_to_bit_it_1_vnu_17_in_0, msg_to_bit_it_1_vnu_17_in_1, msg_to_bit_it_1_vnu_17_in_2, msg_to_bit_it_1_vnu_18_in_0, msg_to_bit_it_1_vnu_18_in_1, msg_to_bit_it_1_vnu_18_in_2, msg_to_bit_it_1_vnu_19_in_0, msg_to_bit_it_1_vnu_19_in_1, msg_to_bit_it_1_vnu_19_in_2, msg_to_bit_it_1_vnu_20_in_0, msg_to_bit_it_1_vnu_20_in_1, msg_to_bit_it_1_vnu_20_in_2, msg_to_bit_it_1_vnu_21_in_0, msg_to_bit_it_1_vnu_21_in_1, msg_to_bit_it_1_vnu_21_in_2, msg_to_bit_it_1_vnu_22_in_0, msg_to_bit_it_1_vnu_22_in_1, msg_to_bit_it_1_vnu_22_in_2, msg_to_bit_it_1_vnu_23_in_0, msg_to_bit_it_1_vnu_23_in_1, msg_to_bit_it_1_vnu_23_in_2, msg_to_bit_it_1_vnu_24_in_0, msg_to_bit_it_1_vnu_24_in_1, msg_to_bit_it_1_vnu_24_in_2, msg_to_bit_it_1_vnu_25_in_0, msg_to_bit_it_1_vnu_25_in_1, msg_to_bit_it_1_vnu_25_in_2, msg_to_bit_it_1_vnu_26_in_0, msg_to_bit_it_1_vnu_26_in_1, msg_to_bit_it_1_vnu_26_in_2, msg_to_bit_it_1_vnu_27_in_0, msg_to_bit_it_1_vnu_27_in_1, msg_to_bit_it_1_vnu_27_in_2, msg_to_bit_it_1_vnu_28_in_0, msg_to_bit_it_1_vnu_28_in_1, msg_to_bit_it_1_vnu_28_in_2, msg_to_bit_it_1_vnu_29_in_0, msg_to_bit_it_1_vnu_29_in_1, msg_to_bit_it_1_vnu_29_in_2, msg_to_bit_it_1_vnu_30_in_0, msg_to_bit_it_1_vnu_30_in_1, msg_to_bit_it_1_vnu_30_in_2, msg_to_bit_it_1_vnu_31_in_0, msg_to_bit_it_1_vnu_31_in_1, msg_to_bit_it_1_vnu_31_in_2, msg_to_bit_it_1_vnu_32_in_0, msg_to_bit_it_1_vnu_32_in_1, msg_to_bit_it_1_vnu_32_in_2, msg_to_bit_it_1_vnu_33_in_0, msg_to_bit_it_1_vnu_33_in_1, msg_to_bit_it_1_vnu_33_in_2, msg_to_bit_it_1_vnu_34_in_0, msg_to_bit_it_1_vnu_34_in_1, msg_to_bit_it_1_vnu_34_in_2, msg_to_bit_it_1_vnu_35_in_0, msg_to_bit_it_1_vnu_35_in_1, msg_to_bit_it_1_vnu_35_in_2, msg_to_bit_it_1_vnu_36_in_0, msg_to_bit_it_1_vnu_36_in_1, msg_to_bit_it_1_vnu_36_in_2, msg_to_bit_it_1_vnu_37_in_0, msg_to_bit_it_1_vnu_37_in_1, msg_to_bit_it_1_vnu_37_in_2, msg_to_bit_it_1_vnu_38_in_0, msg_to_bit_it_1_vnu_38_in_1, msg_to_bit_it_1_vnu_38_in_2, msg_to_bit_it_1_vnu_39_in_0, msg_to_bit_it_1_vnu_39_in_1, msg_to_bit_it_1_vnu_39_in_2, msg_to_bit_it_1_vnu_40_in_0, msg_to_bit_it_1_vnu_40_in_1, msg_to_bit_it_1_vnu_40_in_2, msg_to_bit_it_1_vnu_41_in_0, msg_to_bit_it_1_vnu_41_in_1, msg_to_bit_it_1_vnu_41_in_2, msg_to_bit_it_1_vnu_42_in_0, msg_to_bit_it_1_vnu_42_in_1, msg_to_bit_it_1_vnu_42_in_2, msg_to_bit_it_1_vnu_43_in_0, msg_to_bit_it_1_vnu_43_in_1, msg_to_bit_it_1_vnu_43_in_2, msg_to_bit_it_1_vnu_44_in_0, msg_to_bit_it_1_vnu_44_in_1, msg_to_bit_it_1_vnu_44_in_2, msg_to_bit_it_1_vnu_45_in_0, msg_to_bit_it_1_vnu_45_in_1, msg_to_bit_it_1_vnu_45_in_2, msg_to_bit_it_1_vnu_46_in_0, msg_to_bit_it_1_vnu_46_in_1, msg_to_bit_it_1_vnu_46_in_2, msg_to_bit_it_1_vnu_47_in_0, msg_to_bit_it_1_vnu_47_in_1, msg_to_bit_it_1_vnu_47_in_2, msg_to_bit_it_1_vnu_48_in_0, msg_to_bit_it_1_vnu_48_in_1, msg_to_bit_it_1_vnu_48_in_2, msg_to_bit_it_1_vnu_49_in_0, msg_to_bit_it_1_vnu_49_in_1, msg_to_bit_it_1_vnu_49_in_2, msg_to_bit_it_1_vnu_50_in_0, msg_to_bit_it_1_vnu_50_in_1, msg_to_bit_it_1_vnu_50_in_2, msg_to_bit_it_1_vnu_51_in_0, msg_to_bit_it_1_vnu_51_in_1, msg_to_bit_it_1_vnu_51_in_2, msg_to_bit_it_1_vnu_52_in_0, msg_to_bit_it_1_vnu_52_in_1, msg_to_bit_it_1_vnu_52_in_2, msg_to_bit_it_1_vnu_53_in_0, msg_to_bit_it_1_vnu_53_in_1, msg_to_bit_it_1_vnu_53_in_2, msg_to_bit_it_1_vnu_54_in_0, msg_to_bit_it_1_vnu_54_in_1, msg_to_bit_it_1_vnu_54_in_2, msg_to_bit_it_1_vnu_55_in_0, msg_to_bit_it_1_vnu_55_in_1, msg_to_bit_it_1_vnu_55_in_2, msg_to_bit_it_1_vnu_56_in_0, msg_to_bit_it_1_vnu_56_in_1, msg_to_bit_it_1_vnu_56_in_2, msg_to_bit_it_1_vnu_57_in_0, msg_to_bit_it_1_vnu_57_in_1, msg_to_bit_it_1_vnu_57_in_2, msg_to_bit_it_1_vnu_58_in_0, msg_to_bit_it_1_vnu_58_in_1, msg_to_bit_it_1_vnu_58_in_2, msg_to_bit_it_1_vnu_59_in_0, msg_to_bit_it_1_vnu_59_in_1, msg_to_bit_it_1_vnu_59_in_2, msg_to_bit_it_1_vnu_60_in_0, msg_to_bit_it_1_vnu_60_in_1, msg_to_bit_it_1_vnu_60_in_2, msg_to_bit_it_1_vnu_61_in_0, msg_to_bit_it_1_vnu_61_in_1, msg_to_bit_it_1_vnu_61_in_2, msg_to_bit_it_1_vnu_62_in_0, msg_to_bit_it_1_vnu_62_in_1, msg_to_bit_it_1_vnu_62_in_2, msg_to_bit_it_1_vnu_63_in_0, msg_to_bit_it_1_vnu_63_in_1, msg_to_bit_it_1_vnu_63_in_2, msg_to_bit_it_1_vnu_64_in_0, msg_to_bit_it_1_vnu_64_in_1, msg_to_bit_it_1_vnu_64_in_2, msg_to_bit_it_1_vnu_65_in_0, msg_to_bit_it_1_vnu_65_in_1, msg_to_bit_it_1_vnu_65_in_2, msg_to_bit_it_1_vnu_66_in_0, msg_to_bit_it_1_vnu_66_in_1, msg_to_bit_it_1_vnu_66_in_2, msg_to_bit_it_1_vnu_67_in_0, msg_to_bit_it_1_vnu_67_in_1, msg_to_bit_it_1_vnu_67_in_2, msg_to_bit_it_1_vnu_68_in_0, msg_to_bit_it_1_vnu_68_in_1, msg_to_bit_it_1_vnu_68_in_2, msg_to_bit_it_1_vnu_69_in_0, msg_to_bit_it_1_vnu_69_in_1, msg_to_bit_it_1_vnu_69_in_2, msg_to_bit_it_1_vnu_70_in_0, msg_to_bit_it_1_vnu_70_in_1, msg_to_bit_it_1_vnu_70_in_2, msg_to_bit_it_1_vnu_71_in_0, msg_to_bit_it_1_vnu_71_in_1, msg_to_bit_it_1_vnu_71_in_2, msg_to_bit_it_1_vnu_72_in_0, msg_to_bit_it_1_vnu_72_in_1, msg_to_bit_it_1_vnu_72_in_2, msg_to_bit_it_1_vnu_73_in_0, msg_to_bit_it_1_vnu_73_in_1, msg_to_bit_it_1_vnu_73_in_2, msg_to_bit_it_1_vnu_74_in_0, msg_to_bit_it_1_vnu_74_in_1, msg_to_bit_it_1_vnu_74_in_2, msg_to_bit_it_1_vnu_75_in_0, msg_to_bit_it_1_vnu_75_in_1, msg_to_bit_it_1_vnu_75_in_2, msg_to_bit_it_1_vnu_76_in_0, msg_to_bit_it_1_vnu_76_in_1, msg_to_bit_it_1_vnu_76_in_2, msg_to_bit_it_1_vnu_77_in_0, msg_to_bit_it_1_vnu_77_in_1, msg_to_bit_it_1_vnu_77_in_2, msg_to_bit_it_1_vnu_78_in_0, msg_to_bit_it_1_vnu_78_in_1, msg_to_bit_it_1_vnu_78_in_2, msg_to_bit_it_1_vnu_79_in_0, msg_to_bit_it_1_vnu_79_in_1, msg_to_bit_it_1_vnu_79_in_2, msg_to_bit_it_1_vnu_80_in_0, msg_to_bit_it_1_vnu_80_in_1, msg_to_bit_it_1_vnu_80_in_2, msg_to_bit_it_1_vnu_81_in_0, msg_to_bit_it_1_vnu_81_in_1, msg_to_bit_it_1_vnu_81_in_2, msg_to_bit_it_1_vnu_82_in_0, msg_to_bit_it_1_vnu_82_in_1, msg_to_bit_it_1_vnu_82_in_2, msg_to_bit_it_1_vnu_83_in_0, msg_to_bit_it_1_vnu_83_in_1, msg_to_bit_it_1_vnu_83_in_2, msg_to_bit_it_1_vnu_84_in_0, msg_to_bit_it_1_vnu_84_in_1, msg_to_bit_it_1_vnu_84_in_2, msg_to_bit_it_1_vnu_85_in_0, msg_to_bit_it_1_vnu_85_in_1, msg_to_bit_it_1_vnu_85_in_2, msg_to_bit_it_1_vnu_86_in_0, msg_to_bit_it_1_vnu_86_in_1, msg_to_bit_it_1_vnu_86_in_2, msg_to_bit_it_1_vnu_87_in_0, msg_to_bit_it_1_vnu_87_in_1, msg_to_bit_it_1_vnu_87_in_2, msg_to_bit_it_1_vnu_88_in_0, msg_to_bit_it_1_vnu_88_in_1, msg_to_bit_it_1_vnu_88_in_2, msg_to_bit_it_1_vnu_89_in_0, msg_to_bit_it_1_vnu_89_in_1, msg_to_bit_it_1_vnu_89_in_2, msg_to_bit_it_1_vnu_90_in_0, msg_to_bit_it_1_vnu_90_in_1, msg_to_bit_it_1_vnu_90_in_2, msg_to_bit_it_1_vnu_91_in_0, msg_to_bit_it_1_vnu_91_in_1, msg_to_bit_it_1_vnu_91_in_2, msg_to_bit_it_1_vnu_92_in_0, msg_to_bit_it_1_vnu_92_in_1, msg_to_bit_it_1_vnu_92_in_2, msg_to_bit_it_1_vnu_93_in_0, msg_to_bit_it_1_vnu_93_in_1, msg_to_bit_it_1_vnu_93_in_2, msg_to_bit_it_1_vnu_94_in_0, msg_to_bit_it_1_vnu_94_in_1, msg_to_bit_it_1_vnu_94_in_2, msg_to_bit_it_1_vnu_95_in_0, msg_to_bit_it_1_vnu_95_in_1, msg_to_bit_it_1_vnu_95_in_2, msg_to_bit_it_1_vnu_96_in_0, msg_to_bit_it_1_vnu_96_in_1, msg_to_bit_it_1_vnu_96_in_2, msg_to_bit_it_1_vnu_97_in_0, msg_to_bit_it_1_vnu_97_in_1, msg_to_bit_it_1_vnu_97_in_2, msg_to_bit_it_1_vnu_98_in_0, msg_to_bit_it_1_vnu_98_in_1, msg_to_bit_it_1_vnu_98_in_2, msg_to_bit_it_1_vnu_99_in_0, msg_to_bit_it_1_vnu_99_in_1, msg_to_bit_it_1_vnu_99_in_2, msg_to_bit_it_1_vnu_100_in_0, msg_to_bit_it_1_vnu_100_in_1, msg_to_bit_it_1_vnu_100_in_2, msg_to_bit_it_1_vnu_101_in_0, msg_to_bit_it_1_vnu_101_in_1, msg_to_bit_it_1_vnu_101_in_2, msg_to_bit_it_1_vnu_102_in_0, msg_to_bit_it_1_vnu_102_in_1, msg_to_bit_it_1_vnu_102_in_2, msg_to_bit_it_1_vnu_103_in_0, msg_to_bit_it_1_vnu_103_in_1, msg_to_bit_it_1_vnu_103_in_2, msg_to_bit_it_1_vnu_104_in_0, msg_to_bit_it_1_vnu_104_in_1, msg_to_bit_it_1_vnu_104_in_2, msg_to_bit_it_1_vnu_105_in_0, msg_to_bit_it_1_vnu_105_in_1, msg_to_bit_it_1_vnu_105_in_2, msg_to_bit_it_1_vnu_106_in_0, msg_to_bit_it_1_vnu_106_in_1, msg_to_bit_it_1_vnu_106_in_2, msg_to_bit_it_1_vnu_107_in_0, msg_to_bit_it_1_vnu_107_in_1, msg_to_bit_it_1_vnu_107_in_2, msg_to_bit_it_1_vnu_108_in_0, msg_to_bit_it_1_vnu_108_in_1, msg_to_bit_it_1_vnu_108_in_2, msg_to_bit_it_1_vnu_109_in_0, msg_to_bit_it_1_vnu_109_in_1, msg_to_bit_it_1_vnu_109_in_2, msg_to_bit_it_1_vnu_110_in_0, msg_to_bit_it_1_vnu_110_in_1, msg_to_bit_it_1_vnu_110_in_2, msg_to_bit_it_1_vnu_111_in_0, msg_to_bit_it_1_vnu_111_in_1, msg_to_bit_it_1_vnu_111_in_2, msg_to_bit_it_1_vnu_112_in_0, msg_to_bit_it_1_vnu_112_in_1, msg_to_bit_it_1_vnu_112_in_2, msg_to_bit_it_1_vnu_113_in_0, msg_to_bit_it_1_vnu_113_in_1, msg_to_bit_it_1_vnu_113_in_2, msg_to_bit_it_1_vnu_114_in_0, msg_to_bit_it_1_vnu_114_in_1, msg_to_bit_it_1_vnu_114_in_2, msg_to_bit_it_1_vnu_115_in_0, msg_to_bit_it_1_vnu_115_in_1, msg_to_bit_it_1_vnu_115_in_2, msg_to_bit_it_1_vnu_116_in_0, msg_to_bit_it_1_vnu_116_in_1, msg_to_bit_it_1_vnu_116_in_2, msg_to_bit_it_1_vnu_117_in_0, msg_to_bit_it_1_vnu_117_in_1, msg_to_bit_it_1_vnu_117_in_2, msg_to_bit_it_1_vnu_118_in_0, msg_to_bit_it_1_vnu_118_in_1, msg_to_bit_it_1_vnu_118_in_2, msg_to_bit_it_1_vnu_119_in_0, msg_to_bit_it_1_vnu_119_in_1, msg_to_bit_it_1_vnu_119_in_2, msg_to_bit_it_1_vnu_120_in_0, msg_to_bit_it_1_vnu_120_in_1, msg_to_bit_it_1_vnu_120_in_2, msg_to_bit_it_1_vnu_121_in_0, msg_to_bit_it_1_vnu_121_in_1, msg_to_bit_it_1_vnu_121_in_2, msg_to_bit_it_1_vnu_122_in_0, msg_to_bit_it_1_vnu_122_in_1, msg_to_bit_it_1_vnu_122_in_2, msg_to_bit_it_1_vnu_123_in_0, msg_to_bit_it_1_vnu_123_in_1, msg_to_bit_it_1_vnu_123_in_2, msg_to_bit_it_1_vnu_124_in_0, msg_to_bit_it_1_vnu_124_in_1, msg_to_bit_it_1_vnu_124_in_2, msg_to_bit_it_1_vnu_125_in_0, msg_to_bit_it_1_vnu_125_in_1, msg_to_bit_it_1_vnu_125_in_2, msg_to_bit_it_1_vnu_126_in_0, msg_to_bit_it_1_vnu_126_in_1, msg_to_bit_it_1_vnu_126_in_2, msg_to_bit_it_1_vnu_127_in_0, msg_to_bit_it_1_vnu_127_in_1, msg_to_bit_it_1_vnu_127_in_2, msg_to_bit_it_1_vnu_128_in_0, msg_to_bit_it_1_vnu_128_in_1, msg_to_bit_it_1_vnu_128_in_2, msg_to_bit_it_1_vnu_129_in_0, msg_to_bit_it_1_vnu_129_in_1, msg_to_bit_it_1_vnu_129_in_2, msg_to_bit_it_1_vnu_130_in_0, msg_to_bit_it_1_vnu_130_in_1, msg_to_bit_it_1_vnu_130_in_2, msg_to_bit_it_1_vnu_131_in_0, msg_to_bit_it_1_vnu_131_in_1, msg_to_bit_it_1_vnu_131_in_2, msg_to_bit_it_1_vnu_132_in_0, msg_to_bit_it_1_vnu_132_in_1, msg_to_bit_it_1_vnu_132_in_2, msg_to_bit_it_1_vnu_133_in_0, msg_to_bit_it_1_vnu_133_in_1, msg_to_bit_it_1_vnu_133_in_2, msg_to_bit_it_1_vnu_134_in_0, msg_to_bit_it_1_vnu_134_in_1, msg_to_bit_it_1_vnu_134_in_2, msg_to_bit_it_1_vnu_135_in_0, msg_to_bit_it_1_vnu_135_in_1, msg_to_bit_it_1_vnu_135_in_2, msg_to_bit_it_1_vnu_136_in_0, msg_to_bit_it_1_vnu_136_in_1, msg_to_bit_it_1_vnu_136_in_2, msg_to_bit_it_1_vnu_137_in_0, msg_to_bit_it_1_vnu_137_in_1, msg_to_bit_it_1_vnu_137_in_2, msg_to_bit_it_1_vnu_138_in_0, msg_to_bit_it_1_vnu_138_in_1, msg_to_bit_it_1_vnu_138_in_2, msg_to_bit_it_1_vnu_139_in_0, msg_to_bit_it_1_vnu_139_in_1, msg_to_bit_it_1_vnu_139_in_2, msg_to_bit_it_1_vnu_140_in_0, msg_to_bit_it_1_vnu_140_in_1, msg_to_bit_it_1_vnu_140_in_2, msg_to_bit_it_1_vnu_141_in_0, msg_to_bit_it_1_vnu_141_in_1, msg_to_bit_it_1_vnu_141_in_2, msg_to_bit_it_1_vnu_142_in_0, msg_to_bit_it_1_vnu_142_in_1, msg_to_bit_it_1_vnu_142_in_2, msg_to_bit_it_1_vnu_143_in_0, msg_to_bit_it_1_vnu_143_in_1, msg_to_bit_it_1_vnu_143_in_2, msg_to_bit_it_1_vnu_144_in_0, msg_to_bit_it_1_vnu_144_in_1, msg_to_bit_it_1_vnu_144_in_2, msg_to_bit_it_1_vnu_145_in_0, msg_to_bit_it_1_vnu_145_in_1, msg_to_bit_it_1_vnu_145_in_2, msg_to_bit_it_1_vnu_146_in_0, msg_to_bit_it_1_vnu_146_in_1, msg_to_bit_it_1_vnu_146_in_2, msg_to_bit_it_1_vnu_147_in_0, msg_to_bit_it_1_vnu_147_in_1, msg_to_bit_it_1_vnu_147_in_2, msg_to_bit_it_1_vnu_148_in_0, msg_to_bit_it_1_vnu_148_in_1, msg_to_bit_it_1_vnu_148_in_2, msg_to_bit_it_1_vnu_149_in_0, msg_to_bit_it_1_vnu_149_in_1, msg_to_bit_it_1_vnu_149_in_2, msg_to_bit_it_1_vnu_150_in_0, msg_to_bit_it_1_vnu_150_in_1, msg_to_bit_it_1_vnu_150_in_2, msg_to_bit_it_1_vnu_151_in_0, msg_to_bit_it_1_vnu_151_in_1, msg_to_bit_it_1_vnu_151_in_2, msg_to_bit_it_1_vnu_152_in_0, msg_to_bit_it_1_vnu_152_in_1, msg_to_bit_it_1_vnu_152_in_2, msg_to_bit_it_1_vnu_153_in_0, msg_to_bit_it_1_vnu_153_in_1, msg_to_bit_it_1_vnu_153_in_2, msg_to_bit_it_1_vnu_154_in_0, msg_to_bit_it_1_vnu_154_in_1, msg_to_bit_it_1_vnu_154_in_2, msg_to_bit_it_1_vnu_155_in_0, msg_to_bit_it_1_vnu_155_in_1, msg_to_bit_it_1_vnu_155_in_2, msg_to_bit_it_1_vnu_156_in_0, msg_to_bit_it_1_vnu_156_in_1, msg_to_bit_it_1_vnu_156_in_2, msg_to_bit_it_1_vnu_157_in_0, msg_to_bit_it_1_vnu_157_in_1, msg_to_bit_it_1_vnu_157_in_2, msg_to_bit_it_1_vnu_158_in_0, msg_to_bit_it_1_vnu_158_in_1, msg_to_bit_it_1_vnu_158_in_2, msg_to_bit_it_1_vnu_159_in_0, msg_to_bit_it_1_vnu_159_in_1, msg_to_bit_it_1_vnu_159_in_2, msg_to_bit_it_1_vnu_160_in_0, msg_to_bit_it_1_vnu_160_in_1, msg_to_bit_it_1_vnu_160_in_2, msg_to_bit_it_1_vnu_161_in_0, msg_to_bit_it_1_vnu_161_in_1, msg_to_bit_it_1_vnu_161_in_2, msg_to_bit_it_1_vnu_162_in_0, msg_to_bit_it_1_vnu_162_in_1, msg_to_bit_it_1_vnu_162_in_2, msg_to_bit_it_1_vnu_163_in_0, msg_to_bit_it_1_vnu_163_in_1, msg_to_bit_it_1_vnu_163_in_2, msg_to_bit_it_1_vnu_164_in_0, msg_to_bit_it_1_vnu_164_in_1, msg_to_bit_it_1_vnu_164_in_2, msg_to_bit_it_1_vnu_165_in_0, msg_to_bit_it_1_vnu_165_in_1, msg_to_bit_it_1_vnu_165_in_2, msg_to_bit_it_1_vnu_166_in_0, msg_to_bit_it_1_vnu_166_in_1, msg_to_bit_it_1_vnu_166_in_2, msg_to_bit_it_1_vnu_167_in_0, msg_to_bit_it_1_vnu_167_in_1, msg_to_bit_it_1_vnu_167_in_2, msg_to_bit_it_1_vnu_168_in_0, msg_to_bit_it_1_vnu_168_in_1, msg_to_bit_it_1_vnu_168_in_2, msg_to_bit_it_1_vnu_169_in_0, msg_to_bit_it_1_vnu_169_in_1, msg_to_bit_it_1_vnu_169_in_2, msg_to_bit_it_1_vnu_170_in_0, msg_to_bit_it_1_vnu_170_in_1, msg_to_bit_it_1_vnu_170_in_2, msg_to_bit_it_1_vnu_171_in_0, msg_to_bit_it_1_vnu_171_in_1, msg_to_bit_it_1_vnu_171_in_2, msg_to_bit_it_1_vnu_172_in_0, msg_to_bit_it_1_vnu_172_in_1, msg_to_bit_it_1_vnu_172_in_2, msg_to_bit_it_1_vnu_173_in_0, msg_to_bit_it_1_vnu_173_in_1, msg_to_bit_it_1_vnu_173_in_2, msg_to_bit_it_1_vnu_174_in_0, msg_to_bit_it_1_vnu_174_in_1, msg_to_bit_it_1_vnu_174_in_2, msg_to_bit_it_1_vnu_175_in_0, msg_to_bit_it_1_vnu_175_in_1, msg_to_bit_it_1_vnu_175_in_2, msg_to_bit_it_1_vnu_176_in_0, msg_to_bit_it_1_vnu_176_in_1, msg_to_bit_it_1_vnu_176_in_2, msg_to_bit_it_1_vnu_177_in_0, msg_to_bit_it_1_vnu_177_in_1, msg_to_bit_it_1_vnu_177_in_2, msg_to_bit_it_1_vnu_178_in_0, msg_to_bit_it_1_vnu_178_in_1, msg_to_bit_it_1_vnu_178_in_2, msg_to_bit_it_1_vnu_179_in_0, msg_to_bit_it_1_vnu_179_in_1, msg_to_bit_it_1_vnu_179_in_2, msg_to_bit_it_1_vnu_180_in_0, msg_to_bit_it_1_vnu_180_in_1, msg_to_bit_it_1_vnu_180_in_2, msg_to_bit_it_1_vnu_181_in_0, msg_to_bit_it_1_vnu_181_in_1, msg_to_bit_it_1_vnu_181_in_2, msg_to_bit_it_1_vnu_182_in_0, msg_to_bit_it_1_vnu_182_in_1, msg_to_bit_it_1_vnu_182_in_2, msg_to_bit_it_1_vnu_183_in_0, msg_to_bit_it_1_vnu_183_in_1, msg_to_bit_it_1_vnu_183_in_2, msg_to_bit_it_1_vnu_184_in_0, msg_to_bit_it_1_vnu_184_in_1, msg_to_bit_it_1_vnu_184_in_2, msg_to_bit_it_1_vnu_185_in_0, msg_to_bit_it_1_vnu_185_in_1, msg_to_bit_it_1_vnu_185_in_2, msg_to_bit_it_1_vnu_186_in_0, msg_to_bit_it_1_vnu_186_in_1, msg_to_bit_it_1_vnu_186_in_2, msg_to_bit_it_1_vnu_187_in_0, msg_to_bit_it_1_vnu_187_in_1, msg_to_bit_it_1_vnu_187_in_2, msg_to_bit_it_1_vnu_188_in_0, msg_to_bit_it_1_vnu_188_in_1, msg_to_bit_it_1_vnu_188_in_2, msg_to_bit_it_1_vnu_189_in_0, msg_to_bit_it_1_vnu_189_in_1, msg_to_bit_it_1_vnu_189_in_2, msg_to_bit_it_1_vnu_190_in_0, msg_to_bit_it_1_vnu_190_in_1, msg_to_bit_it_1_vnu_190_in_2, msg_to_bit_it_1_vnu_191_in_0, msg_to_bit_it_1_vnu_191_in_1, msg_to_bit_it_1_vnu_191_in_2, msg_to_bit_it_1_vnu_192_in_0, msg_to_bit_it_1_vnu_192_in_1, msg_to_bit_it_1_vnu_192_in_2, msg_to_bit_it_1_vnu_193_in_0, msg_to_bit_it_1_vnu_193_in_1, msg_to_bit_it_1_vnu_193_in_2, msg_to_bit_it_1_vnu_194_in_0, msg_to_bit_it_1_vnu_194_in_1, msg_to_bit_it_1_vnu_194_in_2, msg_to_bit_it_1_vnu_195_in_0, msg_to_bit_it_1_vnu_195_in_1, msg_to_bit_it_1_vnu_195_in_2, msg_to_bit_it_1_vnu_196_in_0, msg_to_bit_it_1_vnu_196_in_1, msg_to_bit_it_1_vnu_196_in_2, msg_to_bit_it_1_vnu_197_in_0, msg_to_bit_it_1_vnu_197_in_1, msg_to_bit_it_1_vnu_197_in_2, msg_to_bit_it_2_vnu_0_in_0, msg_to_bit_it_2_vnu_0_in_1, msg_to_bit_it_2_vnu_0_in_2, msg_to_bit_it_2_vnu_1_in_0, msg_to_bit_it_2_vnu_1_in_1, msg_to_bit_it_2_vnu_1_in_2, msg_to_bit_it_2_vnu_2_in_0, msg_to_bit_it_2_vnu_2_in_1, msg_to_bit_it_2_vnu_2_in_2, msg_to_bit_it_2_vnu_3_in_0, msg_to_bit_it_2_vnu_3_in_1, msg_to_bit_it_2_vnu_3_in_2, msg_to_bit_it_2_vnu_4_in_0, msg_to_bit_it_2_vnu_4_in_1, msg_to_bit_it_2_vnu_4_in_2, msg_to_bit_it_2_vnu_5_in_0, msg_to_bit_it_2_vnu_5_in_1, msg_to_bit_it_2_vnu_5_in_2, msg_to_bit_it_2_vnu_6_in_0, msg_to_bit_it_2_vnu_6_in_1, msg_to_bit_it_2_vnu_6_in_2, msg_to_bit_it_2_vnu_7_in_0, msg_to_bit_it_2_vnu_7_in_1, msg_to_bit_it_2_vnu_7_in_2, msg_to_bit_it_2_vnu_8_in_0, msg_to_bit_it_2_vnu_8_in_1, msg_to_bit_it_2_vnu_8_in_2, msg_to_bit_it_2_vnu_9_in_0, msg_to_bit_it_2_vnu_9_in_1, msg_to_bit_it_2_vnu_9_in_2, msg_to_bit_it_2_vnu_10_in_0, msg_to_bit_it_2_vnu_10_in_1, msg_to_bit_it_2_vnu_10_in_2, msg_to_bit_it_2_vnu_11_in_0, msg_to_bit_it_2_vnu_11_in_1, msg_to_bit_it_2_vnu_11_in_2, msg_to_bit_it_2_vnu_12_in_0, msg_to_bit_it_2_vnu_12_in_1, msg_to_bit_it_2_vnu_12_in_2, msg_to_bit_it_2_vnu_13_in_0, msg_to_bit_it_2_vnu_13_in_1, msg_to_bit_it_2_vnu_13_in_2, msg_to_bit_it_2_vnu_14_in_0, msg_to_bit_it_2_vnu_14_in_1, msg_to_bit_it_2_vnu_14_in_2, msg_to_bit_it_2_vnu_15_in_0, msg_to_bit_it_2_vnu_15_in_1, msg_to_bit_it_2_vnu_15_in_2, msg_to_bit_it_2_vnu_16_in_0, msg_to_bit_it_2_vnu_16_in_1, msg_to_bit_it_2_vnu_16_in_2, msg_to_bit_it_2_vnu_17_in_0, msg_to_bit_it_2_vnu_17_in_1, msg_to_bit_it_2_vnu_17_in_2, msg_to_bit_it_2_vnu_18_in_0, msg_to_bit_it_2_vnu_18_in_1, msg_to_bit_it_2_vnu_18_in_2, msg_to_bit_it_2_vnu_19_in_0, msg_to_bit_it_2_vnu_19_in_1, msg_to_bit_it_2_vnu_19_in_2, msg_to_bit_it_2_vnu_20_in_0, msg_to_bit_it_2_vnu_20_in_1, msg_to_bit_it_2_vnu_20_in_2, msg_to_bit_it_2_vnu_21_in_0, msg_to_bit_it_2_vnu_21_in_1, msg_to_bit_it_2_vnu_21_in_2, msg_to_bit_it_2_vnu_22_in_0, msg_to_bit_it_2_vnu_22_in_1, msg_to_bit_it_2_vnu_22_in_2, msg_to_bit_it_2_vnu_23_in_0, msg_to_bit_it_2_vnu_23_in_1, msg_to_bit_it_2_vnu_23_in_2, msg_to_bit_it_2_vnu_24_in_0, msg_to_bit_it_2_vnu_24_in_1, msg_to_bit_it_2_vnu_24_in_2, msg_to_bit_it_2_vnu_25_in_0, msg_to_bit_it_2_vnu_25_in_1, msg_to_bit_it_2_vnu_25_in_2, msg_to_bit_it_2_vnu_26_in_0, msg_to_bit_it_2_vnu_26_in_1, msg_to_bit_it_2_vnu_26_in_2, msg_to_bit_it_2_vnu_27_in_0, msg_to_bit_it_2_vnu_27_in_1, msg_to_bit_it_2_vnu_27_in_2, msg_to_bit_it_2_vnu_28_in_0, msg_to_bit_it_2_vnu_28_in_1, msg_to_bit_it_2_vnu_28_in_2, msg_to_bit_it_2_vnu_29_in_0, msg_to_bit_it_2_vnu_29_in_1, msg_to_bit_it_2_vnu_29_in_2, msg_to_bit_it_2_vnu_30_in_0, msg_to_bit_it_2_vnu_30_in_1, msg_to_bit_it_2_vnu_30_in_2, msg_to_bit_it_2_vnu_31_in_0, msg_to_bit_it_2_vnu_31_in_1, msg_to_bit_it_2_vnu_31_in_2, msg_to_bit_it_2_vnu_32_in_0, msg_to_bit_it_2_vnu_32_in_1, msg_to_bit_it_2_vnu_32_in_2, msg_to_bit_it_2_vnu_33_in_0, msg_to_bit_it_2_vnu_33_in_1, msg_to_bit_it_2_vnu_33_in_2, msg_to_bit_it_2_vnu_34_in_0, msg_to_bit_it_2_vnu_34_in_1, msg_to_bit_it_2_vnu_34_in_2, msg_to_bit_it_2_vnu_35_in_0, msg_to_bit_it_2_vnu_35_in_1, msg_to_bit_it_2_vnu_35_in_2, msg_to_bit_it_2_vnu_36_in_0, msg_to_bit_it_2_vnu_36_in_1, msg_to_bit_it_2_vnu_36_in_2, msg_to_bit_it_2_vnu_37_in_0, msg_to_bit_it_2_vnu_37_in_1, msg_to_bit_it_2_vnu_37_in_2, msg_to_bit_it_2_vnu_38_in_0, msg_to_bit_it_2_vnu_38_in_1, msg_to_bit_it_2_vnu_38_in_2, msg_to_bit_it_2_vnu_39_in_0, msg_to_bit_it_2_vnu_39_in_1, msg_to_bit_it_2_vnu_39_in_2, msg_to_bit_it_2_vnu_40_in_0, msg_to_bit_it_2_vnu_40_in_1, msg_to_bit_it_2_vnu_40_in_2, msg_to_bit_it_2_vnu_41_in_0, msg_to_bit_it_2_vnu_41_in_1, msg_to_bit_it_2_vnu_41_in_2, msg_to_bit_it_2_vnu_42_in_0, msg_to_bit_it_2_vnu_42_in_1, msg_to_bit_it_2_vnu_42_in_2, msg_to_bit_it_2_vnu_43_in_0, msg_to_bit_it_2_vnu_43_in_1, msg_to_bit_it_2_vnu_43_in_2, msg_to_bit_it_2_vnu_44_in_0, msg_to_bit_it_2_vnu_44_in_1, msg_to_bit_it_2_vnu_44_in_2, msg_to_bit_it_2_vnu_45_in_0, msg_to_bit_it_2_vnu_45_in_1, msg_to_bit_it_2_vnu_45_in_2, msg_to_bit_it_2_vnu_46_in_0, msg_to_bit_it_2_vnu_46_in_1, msg_to_bit_it_2_vnu_46_in_2, msg_to_bit_it_2_vnu_47_in_0, msg_to_bit_it_2_vnu_47_in_1, msg_to_bit_it_2_vnu_47_in_2, msg_to_bit_it_2_vnu_48_in_0, msg_to_bit_it_2_vnu_48_in_1, msg_to_bit_it_2_vnu_48_in_2, msg_to_bit_it_2_vnu_49_in_0, msg_to_bit_it_2_vnu_49_in_1, msg_to_bit_it_2_vnu_49_in_2, msg_to_bit_it_2_vnu_50_in_0, msg_to_bit_it_2_vnu_50_in_1, msg_to_bit_it_2_vnu_50_in_2, msg_to_bit_it_2_vnu_51_in_0, msg_to_bit_it_2_vnu_51_in_1, msg_to_bit_it_2_vnu_51_in_2, msg_to_bit_it_2_vnu_52_in_0, msg_to_bit_it_2_vnu_52_in_1, msg_to_bit_it_2_vnu_52_in_2, msg_to_bit_it_2_vnu_53_in_0, msg_to_bit_it_2_vnu_53_in_1, msg_to_bit_it_2_vnu_53_in_2, msg_to_bit_it_2_vnu_54_in_0, msg_to_bit_it_2_vnu_54_in_1, msg_to_bit_it_2_vnu_54_in_2, msg_to_bit_it_2_vnu_55_in_0, msg_to_bit_it_2_vnu_55_in_1, msg_to_bit_it_2_vnu_55_in_2, msg_to_bit_it_2_vnu_56_in_0, msg_to_bit_it_2_vnu_56_in_1, msg_to_bit_it_2_vnu_56_in_2, msg_to_bit_it_2_vnu_57_in_0, msg_to_bit_it_2_vnu_57_in_1, msg_to_bit_it_2_vnu_57_in_2, msg_to_bit_it_2_vnu_58_in_0, msg_to_bit_it_2_vnu_58_in_1, msg_to_bit_it_2_vnu_58_in_2, msg_to_bit_it_2_vnu_59_in_0, msg_to_bit_it_2_vnu_59_in_1, msg_to_bit_it_2_vnu_59_in_2, msg_to_bit_it_2_vnu_60_in_0, msg_to_bit_it_2_vnu_60_in_1, msg_to_bit_it_2_vnu_60_in_2, msg_to_bit_it_2_vnu_61_in_0, msg_to_bit_it_2_vnu_61_in_1, msg_to_bit_it_2_vnu_61_in_2, msg_to_bit_it_2_vnu_62_in_0, msg_to_bit_it_2_vnu_62_in_1, msg_to_bit_it_2_vnu_62_in_2, msg_to_bit_it_2_vnu_63_in_0, msg_to_bit_it_2_vnu_63_in_1, msg_to_bit_it_2_vnu_63_in_2, msg_to_bit_it_2_vnu_64_in_0, msg_to_bit_it_2_vnu_64_in_1, msg_to_bit_it_2_vnu_64_in_2, msg_to_bit_it_2_vnu_65_in_0, msg_to_bit_it_2_vnu_65_in_1, msg_to_bit_it_2_vnu_65_in_2, msg_to_bit_it_2_vnu_66_in_0, msg_to_bit_it_2_vnu_66_in_1, msg_to_bit_it_2_vnu_66_in_2, msg_to_bit_it_2_vnu_67_in_0, msg_to_bit_it_2_vnu_67_in_1, msg_to_bit_it_2_vnu_67_in_2, msg_to_bit_it_2_vnu_68_in_0, msg_to_bit_it_2_vnu_68_in_1, msg_to_bit_it_2_vnu_68_in_2, msg_to_bit_it_2_vnu_69_in_0, msg_to_bit_it_2_vnu_69_in_1, msg_to_bit_it_2_vnu_69_in_2, msg_to_bit_it_2_vnu_70_in_0, msg_to_bit_it_2_vnu_70_in_1, msg_to_bit_it_2_vnu_70_in_2, msg_to_bit_it_2_vnu_71_in_0, msg_to_bit_it_2_vnu_71_in_1, msg_to_bit_it_2_vnu_71_in_2, msg_to_bit_it_2_vnu_72_in_0, msg_to_bit_it_2_vnu_72_in_1, msg_to_bit_it_2_vnu_72_in_2, msg_to_bit_it_2_vnu_73_in_0, msg_to_bit_it_2_vnu_73_in_1, msg_to_bit_it_2_vnu_73_in_2, msg_to_bit_it_2_vnu_74_in_0, msg_to_bit_it_2_vnu_74_in_1, msg_to_bit_it_2_vnu_74_in_2, msg_to_bit_it_2_vnu_75_in_0, msg_to_bit_it_2_vnu_75_in_1, msg_to_bit_it_2_vnu_75_in_2, msg_to_bit_it_2_vnu_76_in_0, msg_to_bit_it_2_vnu_76_in_1, msg_to_bit_it_2_vnu_76_in_2, msg_to_bit_it_2_vnu_77_in_0, msg_to_bit_it_2_vnu_77_in_1, msg_to_bit_it_2_vnu_77_in_2, msg_to_bit_it_2_vnu_78_in_0, msg_to_bit_it_2_vnu_78_in_1, msg_to_bit_it_2_vnu_78_in_2, msg_to_bit_it_2_vnu_79_in_0, msg_to_bit_it_2_vnu_79_in_1, msg_to_bit_it_2_vnu_79_in_2, msg_to_bit_it_2_vnu_80_in_0, msg_to_bit_it_2_vnu_80_in_1, msg_to_bit_it_2_vnu_80_in_2, msg_to_bit_it_2_vnu_81_in_0, msg_to_bit_it_2_vnu_81_in_1, msg_to_bit_it_2_vnu_81_in_2, msg_to_bit_it_2_vnu_82_in_0, msg_to_bit_it_2_vnu_82_in_1, msg_to_bit_it_2_vnu_82_in_2, msg_to_bit_it_2_vnu_83_in_0, msg_to_bit_it_2_vnu_83_in_1, msg_to_bit_it_2_vnu_83_in_2, msg_to_bit_it_2_vnu_84_in_0, msg_to_bit_it_2_vnu_84_in_1, msg_to_bit_it_2_vnu_84_in_2, msg_to_bit_it_2_vnu_85_in_0, msg_to_bit_it_2_vnu_85_in_1, msg_to_bit_it_2_vnu_85_in_2, msg_to_bit_it_2_vnu_86_in_0, msg_to_bit_it_2_vnu_86_in_1, msg_to_bit_it_2_vnu_86_in_2, msg_to_bit_it_2_vnu_87_in_0, msg_to_bit_it_2_vnu_87_in_1, msg_to_bit_it_2_vnu_87_in_2, msg_to_bit_it_2_vnu_88_in_0, msg_to_bit_it_2_vnu_88_in_1, msg_to_bit_it_2_vnu_88_in_2, msg_to_bit_it_2_vnu_89_in_0, msg_to_bit_it_2_vnu_89_in_1, msg_to_bit_it_2_vnu_89_in_2, msg_to_bit_it_2_vnu_90_in_0, msg_to_bit_it_2_vnu_90_in_1, msg_to_bit_it_2_vnu_90_in_2, msg_to_bit_it_2_vnu_91_in_0, msg_to_bit_it_2_vnu_91_in_1, msg_to_bit_it_2_vnu_91_in_2, msg_to_bit_it_2_vnu_92_in_0, msg_to_bit_it_2_vnu_92_in_1, msg_to_bit_it_2_vnu_92_in_2, msg_to_bit_it_2_vnu_93_in_0, msg_to_bit_it_2_vnu_93_in_1, msg_to_bit_it_2_vnu_93_in_2, msg_to_bit_it_2_vnu_94_in_0, msg_to_bit_it_2_vnu_94_in_1, msg_to_bit_it_2_vnu_94_in_2, msg_to_bit_it_2_vnu_95_in_0, msg_to_bit_it_2_vnu_95_in_1, msg_to_bit_it_2_vnu_95_in_2, msg_to_bit_it_2_vnu_96_in_0, msg_to_bit_it_2_vnu_96_in_1, msg_to_bit_it_2_vnu_96_in_2, msg_to_bit_it_2_vnu_97_in_0, msg_to_bit_it_2_vnu_97_in_1, msg_to_bit_it_2_vnu_97_in_2, msg_to_bit_it_2_vnu_98_in_0, msg_to_bit_it_2_vnu_98_in_1, msg_to_bit_it_2_vnu_98_in_2, msg_to_bit_it_2_vnu_99_in_0, msg_to_bit_it_2_vnu_99_in_1, msg_to_bit_it_2_vnu_99_in_2, msg_to_bit_it_2_vnu_100_in_0, msg_to_bit_it_2_vnu_100_in_1, msg_to_bit_it_2_vnu_100_in_2, msg_to_bit_it_2_vnu_101_in_0, msg_to_bit_it_2_vnu_101_in_1, msg_to_bit_it_2_vnu_101_in_2, msg_to_bit_it_2_vnu_102_in_0, msg_to_bit_it_2_vnu_102_in_1, msg_to_bit_it_2_vnu_102_in_2, msg_to_bit_it_2_vnu_103_in_0, msg_to_bit_it_2_vnu_103_in_1, msg_to_bit_it_2_vnu_103_in_2, msg_to_bit_it_2_vnu_104_in_0, msg_to_bit_it_2_vnu_104_in_1, msg_to_bit_it_2_vnu_104_in_2, msg_to_bit_it_2_vnu_105_in_0, msg_to_bit_it_2_vnu_105_in_1, msg_to_bit_it_2_vnu_105_in_2, msg_to_bit_it_2_vnu_106_in_0, msg_to_bit_it_2_vnu_106_in_1, msg_to_bit_it_2_vnu_106_in_2, msg_to_bit_it_2_vnu_107_in_0, msg_to_bit_it_2_vnu_107_in_1, msg_to_bit_it_2_vnu_107_in_2, msg_to_bit_it_2_vnu_108_in_0, msg_to_bit_it_2_vnu_108_in_1, msg_to_bit_it_2_vnu_108_in_2, msg_to_bit_it_2_vnu_109_in_0, msg_to_bit_it_2_vnu_109_in_1, msg_to_bit_it_2_vnu_109_in_2, msg_to_bit_it_2_vnu_110_in_0, msg_to_bit_it_2_vnu_110_in_1, msg_to_bit_it_2_vnu_110_in_2, msg_to_bit_it_2_vnu_111_in_0, msg_to_bit_it_2_vnu_111_in_1, msg_to_bit_it_2_vnu_111_in_2, msg_to_bit_it_2_vnu_112_in_0, msg_to_bit_it_2_vnu_112_in_1, msg_to_bit_it_2_vnu_112_in_2, msg_to_bit_it_2_vnu_113_in_0, msg_to_bit_it_2_vnu_113_in_1, msg_to_bit_it_2_vnu_113_in_2, msg_to_bit_it_2_vnu_114_in_0, msg_to_bit_it_2_vnu_114_in_1, msg_to_bit_it_2_vnu_114_in_2, msg_to_bit_it_2_vnu_115_in_0, msg_to_bit_it_2_vnu_115_in_1, msg_to_bit_it_2_vnu_115_in_2, msg_to_bit_it_2_vnu_116_in_0, msg_to_bit_it_2_vnu_116_in_1, msg_to_bit_it_2_vnu_116_in_2, msg_to_bit_it_2_vnu_117_in_0, msg_to_bit_it_2_vnu_117_in_1, msg_to_bit_it_2_vnu_117_in_2, msg_to_bit_it_2_vnu_118_in_0, msg_to_bit_it_2_vnu_118_in_1, msg_to_bit_it_2_vnu_118_in_2, msg_to_bit_it_2_vnu_119_in_0, msg_to_bit_it_2_vnu_119_in_1, msg_to_bit_it_2_vnu_119_in_2, msg_to_bit_it_2_vnu_120_in_0, msg_to_bit_it_2_vnu_120_in_1, msg_to_bit_it_2_vnu_120_in_2, msg_to_bit_it_2_vnu_121_in_0, msg_to_bit_it_2_vnu_121_in_1, msg_to_bit_it_2_vnu_121_in_2, msg_to_bit_it_2_vnu_122_in_0, msg_to_bit_it_2_vnu_122_in_1, msg_to_bit_it_2_vnu_122_in_2, msg_to_bit_it_2_vnu_123_in_0, msg_to_bit_it_2_vnu_123_in_1, msg_to_bit_it_2_vnu_123_in_2, msg_to_bit_it_2_vnu_124_in_0, msg_to_bit_it_2_vnu_124_in_1, msg_to_bit_it_2_vnu_124_in_2, msg_to_bit_it_2_vnu_125_in_0, msg_to_bit_it_2_vnu_125_in_1, msg_to_bit_it_2_vnu_125_in_2, msg_to_bit_it_2_vnu_126_in_0, msg_to_bit_it_2_vnu_126_in_1, msg_to_bit_it_2_vnu_126_in_2, msg_to_bit_it_2_vnu_127_in_0, msg_to_bit_it_2_vnu_127_in_1, msg_to_bit_it_2_vnu_127_in_2, msg_to_bit_it_2_vnu_128_in_0, msg_to_bit_it_2_vnu_128_in_1, msg_to_bit_it_2_vnu_128_in_2, msg_to_bit_it_2_vnu_129_in_0, msg_to_bit_it_2_vnu_129_in_1, msg_to_bit_it_2_vnu_129_in_2, msg_to_bit_it_2_vnu_130_in_0, msg_to_bit_it_2_vnu_130_in_1, msg_to_bit_it_2_vnu_130_in_2, msg_to_bit_it_2_vnu_131_in_0, msg_to_bit_it_2_vnu_131_in_1, msg_to_bit_it_2_vnu_131_in_2, msg_to_bit_it_2_vnu_132_in_0, msg_to_bit_it_2_vnu_132_in_1, msg_to_bit_it_2_vnu_132_in_2, msg_to_bit_it_2_vnu_133_in_0, msg_to_bit_it_2_vnu_133_in_1, msg_to_bit_it_2_vnu_133_in_2, msg_to_bit_it_2_vnu_134_in_0, msg_to_bit_it_2_vnu_134_in_1, msg_to_bit_it_2_vnu_134_in_2, msg_to_bit_it_2_vnu_135_in_0, msg_to_bit_it_2_vnu_135_in_1, msg_to_bit_it_2_vnu_135_in_2, msg_to_bit_it_2_vnu_136_in_0, msg_to_bit_it_2_vnu_136_in_1, msg_to_bit_it_2_vnu_136_in_2, msg_to_bit_it_2_vnu_137_in_0, msg_to_bit_it_2_vnu_137_in_1, msg_to_bit_it_2_vnu_137_in_2, msg_to_bit_it_2_vnu_138_in_0, msg_to_bit_it_2_vnu_138_in_1, msg_to_bit_it_2_vnu_138_in_2, msg_to_bit_it_2_vnu_139_in_0, msg_to_bit_it_2_vnu_139_in_1, msg_to_bit_it_2_vnu_139_in_2, msg_to_bit_it_2_vnu_140_in_0, msg_to_bit_it_2_vnu_140_in_1, msg_to_bit_it_2_vnu_140_in_2, msg_to_bit_it_2_vnu_141_in_0, msg_to_bit_it_2_vnu_141_in_1, msg_to_bit_it_2_vnu_141_in_2, msg_to_bit_it_2_vnu_142_in_0, msg_to_bit_it_2_vnu_142_in_1, msg_to_bit_it_2_vnu_142_in_2, msg_to_bit_it_2_vnu_143_in_0, msg_to_bit_it_2_vnu_143_in_1, msg_to_bit_it_2_vnu_143_in_2, msg_to_bit_it_2_vnu_144_in_0, msg_to_bit_it_2_vnu_144_in_1, msg_to_bit_it_2_vnu_144_in_2, msg_to_bit_it_2_vnu_145_in_0, msg_to_bit_it_2_vnu_145_in_1, msg_to_bit_it_2_vnu_145_in_2, msg_to_bit_it_2_vnu_146_in_0, msg_to_bit_it_2_vnu_146_in_1, msg_to_bit_it_2_vnu_146_in_2, msg_to_bit_it_2_vnu_147_in_0, msg_to_bit_it_2_vnu_147_in_1, msg_to_bit_it_2_vnu_147_in_2, msg_to_bit_it_2_vnu_148_in_0, msg_to_bit_it_2_vnu_148_in_1, msg_to_bit_it_2_vnu_148_in_2, msg_to_bit_it_2_vnu_149_in_0, msg_to_bit_it_2_vnu_149_in_1, msg_to_bit_it_2_vnu_149_in_2, msg_to_bit_it_2_vnu_150_in_0, msg_to_bit_it_2_vnu_150_in_1, msg_to_bit_it_2_vnu_150_in_2, msg_to_bit_it_2_vnu_151_in_0, msg_to_bit_it_2_vnu_151_in_1, msg_to_bit_it_2_vnu_151_in_2, msg_to_bit_it_2_vnu_152_in_0, msg_to_bit_it_2_vnu_152_in_1, msg_to_bit_it_2_vnu_152_in_2, msg_to_bit_it_2_vnu_153_in_0, msg_to_bit_it_2_vnu_153_in_1, msg_to_bit_it_2_vnu_153_in_2, msg_to_bit_it_2_vnu_154_in_0, msg_to_bit_it_2_vnu_154_in_1, msg_to_bit_it_2_vnu_154_in_2, msg_to_bit_it_2_vnu_155_in_0, msg_to_bit_it_2_vnu_155_in_1, msg_to_bit_it_2_vnu_155_in_2, msg_to_bit_it_2_vnu_156_in_0, msg_to_bit_it_2_vnu_156_in_1, msg_to_bit_it_2_vnu_156_in_2, msg_to_bit_it_2_vnu_157_in_0, msg_to_bit_it_2_vnu_157_in_1, msg_to_bit_it_2_vnu_157_in_2, msg_to_bit_it_2_vnu_158_in_0, msg_to_bit_it_2_vnu_158_in_1, msg_to_bit_it_2_vnu_158_in_2, msg_to_bit_it_2_vnu_159_in_0, msg_to_bit_it_2_vnu_159_in_1, msg_to_bit_it_2_vnu_159_in_2, msg_to_bit_it_2_vnu_160_in_0, msg_to_bit_it_2_vnu_160_in_1, msg_to_bit_it_2_vnu_160_in_2, msg_to_bit_it_2_vnu_161_in_0, msg_to_bit_it_2_vnu_161_in_1, msg_to_bit_it_2_vnu_161_in_2, msg_to_bit_it_2_vnu_162_in_0, msg_to_bit_it_2_vnu_162_in_1, msg_to_bit_it_2_vnu_162_in_2, msg_to_bit_it_2_vnu_163_in_0, msg_to_bit_it_2_vnu_163_in_1, msg_to_bit_it_2_vnu_163_in_2, msg_to_bit_it_2_vnu_164_in_0, msg_to_bit_it_2_vnu_164_in_1, msg_to_bit_it_2_vnu_164_in_2, msg_to_bit_it_2_vnu_165_in_0, msg_to_bit_it_2_vnu_165_in_1, msg_to_bit_it_2_vnu_165_in_2, msg_to_bit_it_2_vnu_166_in_0, msg_to_bit_it_2_vnu_166_in_1, msg_to_bit_it_2_vnu_166_in_2, msg_to_bit_it_2_vnu_167_in_0, msg_to_bit_it_2_vnu_167_in_1, msg_to_bit_it_2_vnu_167_in_2, msg_to_bit_it_2_vnu_168_in_0, msg_to_bit_it_2_vnu_168_in_1, msg_to_bit_it_2_vnu_168_in_2, msg_to_bit_it_2_vnu_169_in_0, msg_to_bit_it_2_vnu_169_in_1, msg_to_bit_it_2_vnu_169_in_2, msg_to_bit_it_2_vnu_170_in_0, msg_to_bit_it_2_vnu_170_in_1, msg_to_bit_it_2_vnu_170_in_2, msg_to_bit_it_2_vnu_171_in_0, msg_to_bit_it_2_vnu_171_in_1, msg_to_bit_it_2_vnu_171_in_2, msg_to_bit_it_2_vnu_172_in_0, msg_to_bit_it_2_vnu_172_in_1, msg_to_bit_it_2_vnu_172_in_2, msg_to_bit_it_2_vnu_173_in_0, msg_to_bit_it_2_vnu_173_in_1, msg_to_bit_it_2_vnu_173_in_2, msg_to_bit_it_2_vnu_174_in_0, msg_to_bit_it_2_vnu_174_in_1, msg_to_bit_it_2_vnu_174_in_2, msg_to_bit_it_2_vnu_175_in_0, msg_to_bit_it_2_vnu_175_in_1, msg_to_bit_it_2_vnu_175_in_2, msg_to_bit_it_2_vnu_176_in_0, msg_to_bit_it_2_vnu_176_in_1, msg_to_bit_it_2_vnu_176_in_2, msg_to_bit_it_2_vnu_177_in_0, msg_to_bit_it_2_vnu_177_in_1, msg_to_bit_it_2_vnu_177_in_2, msg_to_bit_it_2_vnu_178_in_0, msg_to_bit_it_2_vnu_178_in_1, msg_to_bit_it_2_vnu_178_in_2, msg_to_bit_it_2_vnu_179_in_0, msg_to_bit_it_2_vnu_179_in_1, msg_to_bit_it_2_vnu_179_in_2, msg_to_bit_it_2_vnu_180_in_0, msg_to_bit_it_2_vnu_180_in_1, msg_to_bit_it_2_vnu_180_in_2, msg_to_bit_it_2_vnu_181_in_0, msg_to_bit_it_2_vnu_181_in_1, msg_to_bit_it_2_vnu_181_in_2, msg_to_bit_it_2_vnu_182_in_0, msg_to_bit_it_2_vnu_182_in_1, msg_to_bit_it_2_vnu_182_in_2, msg_to_bit_it_2_vnu_183_in_0, msg_to_bit_it_2_vnu_183_in_1, msg_to_bit_it_2_vnu_183_in_2, msg_to_bit_it_2_vnu_184_in_0, msg_to_bit_it_2_vnu_184_in_1, msg_to_bit_it_2_vnu_184_in_2, msg_to_bit_it_2_vnu_185_in_0, msg_to_bit_it_2_vnu_185_in_1, msg_to_bit_it_2_vnu_185_in_2, msg_to_bit_it_2_vnu_186_in_0, msg_to_bit_it_2_vnu_186_in_1, msg_to_bit_it_2_vnu_186_in_2, msg_to_bit_it_2_vnu_187_in_0, msg_to_bit_it_2_vnu_187_in_1, msg_to_bit_it_2_vnu_187_in_2, msg_to_bit_it_2_vnu_188_in_0, msg_to_bit_it_2_vnu_188_in_1, msg_to_bit_it_2_vnu_188_in_2, msg_to_bit_it_2_vnu_189_in_0, msg_to_bit_it_2_vnu_189_in_1, msg_to_bit_it_2_vnu_189_in_2, msg_to_bit_it_2_vnu_190_in_0, msg_to_bit_it_2_vnu_190_in_1, msg_to_bit_it_2_vnu_190_in_2, msg_to_bit_it_2_vnu_191_in_0, msg_to_bit_it_2_vnu_191_in_1, msg_to_bit_it_2_vnu_191_in_2, msg_to_bit_it_2_vnu_192_in_0, msg_to_bit_it_2_vnu_192_in_1, msg_to_bit_it_2_vnu_192_in_2, msg_to_bit_it_2_vnu_193_in_0, msg_to_bit_it_2_vnu_193_in_1, msg_to_bit_it_2_vnu_193_in_2, msg_to_bit_it_2_vnu_194_in_0, msg_to_bit_it_2_vnu_194_in_1, msg_to_bit_it_2_vnu_194_in_2, msg_to_bit_it_2_vnu_195_in_0, msg_to_bit_it_2_vnu_195_in_1, msg_to_bit_it_2_vnu_195_in_2, msg_to_bit_it_2_vnu_196_in_0, msg_to_bit_it_2_vnu_196_in_1, msg_to_bit_it_2_vnu_196_in_2, msg_to_bit_it_2_vnu_197_in_0, msg_to_bit_it_2_vnu_197_in_1, msg_to_bit_it_2_vnu_197_in_2, msg_to_bit_it_3_vnu_0_in_0, msg_to_bit_it_3_vnu_0_in_1, msg_to_bit_it_3_vnu_0_in_2, msg_to_bit_it_3_vnu_1_in_0, msg_to_bit_it_3_vnu_1_in_1, msg_to_bit_it_3_vnu_1_in_2, msg_to_bit_it_3_vnu_2_in_0, msg_to_bit_it_3_vnu_2_in_1, msg_to_bit_it_3_vnu_2_in_2, msg_to_bit_it_3_vnu_3_in_0, msg_to_bit_it_3_vnu_3_in_1, msg_to_bit_it_3_vnu_3_in_2, msg_to_bit_it_3_vnu_4_in_0, msg_to_bit_it_3_vnu_4_in_1, msg_to_bit_it_3_vnu_4_in_2, msg_to_bit_it_3_vnu_5_in_0, msg_to_bit_it_3_vnu_5_in_1, msg_to_bit_it_3_vnu_5_in_2, msg_to_bit_it_3_vnu_6_in_0, msg_to_bit_it_3_vnu_6_in_1, msg_to_bit_it_3_vnu_6_in_2, msg_to_bit_it_3_vnu_7_in_0, msg_to_bit_it_3_vnu_7_in_1, msg_to_bit_it_3_vnu_7_in_2, msg_to_bit_it_3_vnu_8_in_0, msg_to_bit_it_3_vnu_8_in_1, msg_to_bit_it_3_vnu_8_in_2, msg_to_bit_it_3_vnu_9_in_0, msg_to_bit_it_3_vnu_9_in_1, msg_to_bit_it_3_vnu_9_in_2, msg_to_bit_it_3_vnu_10_in_0, msg_to_bit_it_3_vnu_10_in_1, msg_to_bit_it_3_vnu_10_in_2, msg_to_bit_it_3_vnu_11_in_0, msg_to_bit_it_3_vnu_11_in_1, msg_to_bit_it_3_vnu_11_in_2, msg_to_bit_it_3_vnu_12_in_0, msg_to_bit_it_3_vnu_12_in_1, msg_to_bit_it_3_vnu_12_in_2, msg_to_bit_it_3_vnu_13_in_0, msg_to_bit_it_3_vnu_13_in_1, msg_to_bit_it_3_vnu_13_in_2, msg_to_bit_it_3_vnu_14_in_0, msg_to_bit_it_3_vnu_14_in_1, msg_to_bit_it_3_vnu_14_in_2, msg_to_bit_it_3_vnu_15_in_0, msg_to_bit_it_3_vnu_15_in_1, msg_to_bit_it_3_vnu_15_in_2, msg_to_bit_it_3_vnu_16_in_0, msg_to_bit_it_3_vnu_16_in_1, msg_to_bit_it_3_vnu_16_in_2, msg_to_bit_it_3_vnu_17_in_0, msg_to_bit_it_3_vnu_17_in_1, msg_to_bit_it_3_vnu_17_in_2, msg_to_bit_it_3_vnu_18_in_0, msg_to_bit_it_3_vnu_18_in_1, msg_to_bit_it_3_vnu_18_in_2, msg_to_bit_it_3_vnu_19_in_0, msg_to_bit_it_3_vnu_19_in_1, msg_to_bit_it_3_vnu_19_in_2, msg_to_bit_it_3_vnu_20_in_0, msg_to_bit_it_3_vnu_20_in_1, msg_to_bit_it_3_vnu_20_in_2, msg_to_bit_it_3_vnu_21_in_0, msg_to_bit_it_3_vnu_21_in_1, msg_to_bit_it_3_vnu_21_in_2, msg_to_bit_it_3_vnu_22_in_0, msg_to_bit_it_3_vnu_22_in_1, msg_to_bit_it_3_vnu_22_in_2, msg_to_bit_it_3_vnu_23_in_0, msg_to_bit_it_3_vnu_23_in_1, msg_to_bit_it_3_vnu_23_in_2, msg_to_bit_it_3_vnu_24_in_0, msg_to_bit_it_3_vnu_24_in_1, msg_to_bit_it_3_vnu_24_in_2, msg_to_bit_it_3_vnu_25_in_0, msg_to_bit_it_3_vnu_25_in_1, msg_to_bit_it_3_vnu_25_in_2, msg_to_bit_it_3_vnu_26_in_0, msg_to_bit_it_3_vnu_26_in_1, msg_to_bit_it_3_vnu_26_in_2, msg_to_bit_it_3_vnu_27_in_0, msg_to_bit_it_3_vnu_27_in_1, msg_to_bit_it_3_vnu_27_in_2, msg_to_bit_it_3_vnu_28_in_0, msg_to_bit_it_3_vnu_28_in_1, msg_to_bit_it_3_vnu_28_in_2, msg_to_bit_it_3_vnu_29_in_0, msg_to_bit_it_3_vnu_29_in_1, msg_to_bit_it_3_vnu_29_in_2, msg_to_bit_it_3_vnu_30_in_0, msg_to_bit_it_3_vnu_30_in_1, msg_to_bit_it_3_vnu_30_in_2, msg_to_bit_it_3_vnu_31_in_0, msg_to_bit_it_3_vnu_31_in_1, msg_to_bit_it_3_vnu_31_in_2, msg_to_bit_it_3_vnu_32_in_0, msg_to_bit_it_3_vnu_32_in_1, msg_to_bit_it_3_vnu_32_in_2, msg_to_bit_it_3_vnu_33_in_0, msg_to_bit_it_3_vnu_33_in_1, msg_to_bit_it_3_vnu_33_in_2, msg_to_bit_it_3_vnu_34_in_0, msg_to_bit_it_3_vnu_34_in_1, msg_to_bit_it_3_vnu_34_in_2, msg_to_bit_it_3_vnu_35_in_0, msg_to_bit_it_3_vnu_35_in_1, msg_to_bit_it_3_vnu_35_in_2, msg_to_bit_it_3_vnu_36_in_0, msg_to_bit_it_3_vnu_36_in_1, msg_to_bit_it_3_vnu_36_in_2, msg_to_bit_it_3_vnu_37_in_0, msg_to_bit_it_3_vnu_37_in_1, msg_to_bit_it_3_vnu_37_in_2, msg_to_bit_it_3_vnu_38_in_0, msg_to_bit_it_3_vnu_38_in_1, msg_to_bit_it_3_vnu_38_in_2, msg_to_bit_it_3_vnu_39_in_0, msg_to_bit_it_3_vnu_39_in_1, msg_to_bit_it_3_vnu_39_in_2, msg_to_bit_it_3_vnu_40_in_0, msg_to_bit_it_3_vnu_40_in_1, msg_to_bit_it_3_vnu_40_in_2, msg_to_bit_it_3_vnu_41_in_0, msg_to_bit_it_3_vnu_41_in_1, msg_to_bit_it_3_vnu_41_in_2, msg_to_bit_it_3_vnu_42_in_0, msg_to_bit_it_3_vnu_42_in_1, msg_to_bit_it_3_vnu_42_in_2, msg_to_bit_it_3_vnu_43_in_0, msg_to_bit_it_3_vnu_43_in_1, msg_to_bit_it_3_vnu_43_in_2, msg_to_bit_it_3_vnu_44_in_0, msg_to_bit_it_3_vnu_44_in_1, msg_to_bit_it_3_vnu_44_in_2, msg_to_bit_it_3_vnu_45_in_0, msg_to_bit_it_3_vnu_45_in_1, msg_to_bit_it_3_vnu_45_in_2, msg_to_bit_it_3_vnu_46_in_0, msg_to_bit_it_3_vnu_46_in_1, msg_to_bit_it_3_vnu_46_in_2, msg_to_bit_it_3_vnu_47_in_0, msg_to_bit_it_3_vnu_47_in_1, msg_to_bit_it_3_vnu_47_in_2, msg_to_bit_it_3_vnu_48_in_0, msg_to_bit_it_3_vnu_48_in_1, msg_to_bit_it_3_vnu_48_in_2, msg_to_bit_it_3_vnu_49_in_0, msg_to_bit_it_3_vnu_49_in_1, msg_to_bit_it_3_vnu_49_in_2, msg_to_bit_it_3_vnu_50_in_0, msg_to_bit_it_3_vnu_50_in_1, msg_to_bit_it_3_vnu_50_in_2, msg_to_bit_it_3_vnu_51_in_0, msg_to_bit_it_3_vnu_51_in_1, msg_to_bit_it_3_vnu_51_in_2, msg_to_bit_it_3_vnu_52_in_0, msg_to_bit_it_3_vnu_52_in_1, msg_to_bit_it_3_vnu_52_in_2, msg_to_bit_it_3_vnu_53_in_0, msg_to_bit_it_3_vnu_53_in_1, msg_to_bit_it_3_vnu_53_in_2, msg_to_bit_it_3_vnu_54_in_0, msg_to_bit_it_3_vnu_54_in_1, msg_to_bit_it_3_vnu_54_in_2, msg_to_bit_it_3_vnu_55_in_0, msg_to_bit_it_3_vnu_55_in_1, msg_to_bit_it_3_vnu_55_in_2, msg_to_bit_it_3_vnu_56_in_0, msg_to_bit_it_3_vnu_56_in_1, msg_to_bit_it_3_vnu_56_in_2, msg_to_bit_it_3_vnu_57_in_0, msg_to_bit_it_3_vnu_57_in_1, msg_to_bit_it_3_vnu_57_in_2, msg_to_bit_it_3_vnu_58_in_0, msg_to_bit_it_3_vnu_58_in_1, msg_to_bit_it_3_vnu_58_in_2, msg_to_bit_it_3_vnu_59_in_0, msg_to_bit_it_3_vnu_59_in_1, msg_to_bit_it_3_vnu_59_in_2, msg_to_bit_it_3_vnu_60_in_0, msg_to_bit_it_3_vnu_60_in_1, msg_to_bit_it_3_vnu_60_in_2, msg_to_bit_it_3_vnu_61_in_0, msg_to_bit_it_3_vnu_61_in_1, msg_to_bit_it_3_vnu_61_in_2, msg_to_bit_it_3_vnu_62_in_0, msg_to_bit_it_3_vnu_62_in_1, msg_to_bit_it_3_vnu_62_in_2, msg_to_bit_it_3_vnu_63_in_0, msg_to_bit_it_3_vnu_63_in_1, msg_to_bit_it_3_vnu_63_in_2, msg_to_bit_it_3_vnu_64_in_0, msg_to_bit_it_3_vnu_64_in_1, msg_to_bit_it_3_vnu_64_in_2, msg_to_bit_it_3_vnu_65_in_0, msg_to_bit_it_3_vnu_65_in_1, msg_to_bit_it_3_vnu_65_in_2, msg_to_bit_it_3_vnu_66_in_0, msg_to_bit_it_3_vnu_66_in_1, msg_to_bit_it_3_vnu_66_in_2, msg_to_bit_it_3_vnu_67_in_0, msg_to_bit_it_3_vnu_67_in_1, msg_to_bit_it_3_vnu_67_in_2, msg_to_bit_it_3_vnu_68_in_0, msg_to_bit_it_3_vnu_68_in_1, msg_to_bit_it_3_vnu_68_in_2, msg_to_bit_it_3_vnu_69_in_0, msg_to_bit_it_3_vnu_69_in_1, msg_to_bit_it_3_vnu_69_in_2, msg_to_bit_it_3_vnu_70_in_0, msg_to_bit_it_3_vnu_70_in_1, msg_to_bit_it_3_vnu_70_in_2, msg_to_bit_it_3_vnu_71_in_0, msg_to_bit_it_3_vnu_71_in_1, msg_to_bit_it_3_vnu_71_in_2, msg_to_bit_it_3_vnu_72_in_0, msg_to_bit_it_3_vnu_72_in_1, msg_to_bit_it_3_vnu_72_in_2, msg_to_bit_it_3_vnu_73_in_0, msg_to_bit_it_3_vnu_73_in_1, msg_to_bit_it_3_vnu_73_in_2, msg_to_bit_it_3_vnu_74_in_0, msg_to_bit_it_3_vnu_74_in_1, msg_to_bit_it_3_vnu_74_in_2, msg_to_bit_it_3_vnu_75_in_0, msg_to_bit_it_3_vnu_75_in_1, msg_to_bit_it_3_vnu_75_in_2, msg_to_bit_it_3_vnu_76_in_0, msg_to_bit_it_3_vnu_76_in_1, msg_to_bit_it_3_vnu_76_in_2, msg_to_bit_it_3_vnu_77_in_0, msg_to_bit_it_3_vnu_77_in_1, msg_to_bit_it_3_vnu_77_in_2, msg_to_bit_it_3_vnu_78_in_0, msg_to_bit_it_3_vnu_78_in_1, msg_to_bit_it_3_vnu_78_in_2, msg_to_bit_it_3_vnu_79_in_0, msg_to_bit_it_3_vnu_79_in_1, msg_to_bit_it_3_vnu_79_in_2, msg_to_bit_it_3_vnu_80_in_0, msg_to_bit_it_3_vnu_80_in_1, msg_to_bit_it_3_vnu_80_in_2, msg_to_bit_it_3_vnu_81_in_0, msg_to_bit_it_3_vnu_81_in_1, msg_to_bit_it_3_vnu_81_in_2, msg_to_bit_it_3_vnu_82_in_0, msg_to_bit_it_3_vnu_82_in_1, msg_to_bit_it_3_vnu_82_in_2, msg_to_bit_it_3_vnu_83_in_0, msg_to_bit_it_3_vnu_83_in_1, msg_to_bit_it_3_vnu_83_in_2, msg_to_bit_it_3_vnu_84_in_0, msg_to_bit_it_3_vnu_84_in_1, msg_to_bit_it_3_vnu_84_in_2, msg_to_bit_it_3_vnu_85_in_0, msg_to_bit_it_3_vnu_85_in_1, msg_to_bit_it_3_vnu_85_in_2, msg_to_bit_it_3_vnu_86_in_0, msg_to_bit_it_3_vnu_86_in_1, msg_to_bit_it_3_vnu_86_in_2, msg_to_bit_it_3_vnu_87_in_0, msg_to_bit_it_3_vnu_87_in_1, msg_to_bit_it_3_vnu_87_in_2, msg_to_bit_it_3_vnu_88_in_0, msg_to_bit_it_3_vnu_88_in_1, msg_to_bit_it_3_vnu_88_in_2, msg_to_bit_it_3_vnu_89_in_0, msg_to_bit_it_3_vnu_89_in_1, msg_to_bit_it_3_vnu_89_in_2, msg_to_bit_it_3_vnu_90_in_0, msg_to_bit_it_3_vnu_90_in_1, msg_to_bit_it_3_vnu_90_in_2, msg_to_bit_it_3_vnu_91_in_0, msg_to_bit_it_3_vnu_91_in_1, msg_to_bit_it_3_vnu_91_in_2, msg_to_bit_it_3_vnu_92_in_0, msg_to_bit_it_3_vnu_92_in_1, msg_to_bit_it_3_vnu_92_in_2, msg_to_bit_it_3_vnu_93_in_0, msg_to_bit_it_3_vnu_93_in_1, msg_to_bit_it_3_vnu_93_in_2, msg_to_bit_it_3_vnu_94_in_0, msg_to_bit_it_3_vnu_94_in_1, msg_to_bit_it_3_vnu_94_in_2, msg_to_bit_it_3_vnu_95_in_0, msg_to_bit_it_3_vnu_95_in_1, msg_to_bit_it_3_vnu_95_in_2, msg_to_bit_it_3_vnu_96_in_0, msg_to_bit_it_3_vnu_96_in_1, msg_to_bit_it_3_vnu_96_in_2, msg_to_bit_it_3_vnu_97_in_0, msg_to_bit_it_3_vnu_97_in_1, msg_to_bit_it_3_vnu_97_in_2, msg_to_bit_it_3_vnu_98_in_0, msg_to_bit_it_3_vnu_98_in_1, msg_to_bit_it_3_vnu_98_in_2, msg_to_bit_it_3_vnu_99_in_0, msg_to_bit_it_3_vnu_99_in_1, msg_to_bit_it_3_vnu_99_in_2, msg_to_bit_it_3_vnu_100_in_0, msg_to_bit_it_3_vnu_100_in_1, msg_to_bit_it_3_vnu_100_in_2, msg_to_bit_it_3_vnu_101_in_0, msg_to_bit_it_3_vnu_101_in_1, msg_to_bit_it_3_vnu_101_in_2, msg_to_bit_it_3_vnu_102_in_0, msg_to_bit_it_3_vnu_102_in_1, msg_to_bit_it_3_vnu_102_in_2, msg_to_bit_it_3_vnu_103_in_0, msg_to_bit_it_3_vnu_103_in_1, msg_to_bit_it_3_vnu_103_in_2, msg_to_bit_it_3_vnu_104_in_0, msg_to_bit_it_3_vnu_104_in_1, msg_to_bit_it_3_vnu_104_in_2, msg_to_bit_it_3_vnu_105_in_0, msg_to_bit_it_3_vnu_105_in_1, msg_to_bit_it_3_vnu_105_in_2, msg_to_bit_it_3_vnu_106_in_0, msg_to_bit_it_3_vnu_106_in_1, msg_to_bit_it_3_vnu_106_in_2, msg_to_bit_it_3_vnu_107_in_0, msg_to_bit_it_3_vnu_107_in_1, msg_to_bit_it_3_vnu_107_in_2, msg_to_bit_it_3_vnu_108_in_0, msg_to_bit_it_3_vnu_108_in_1, msg_to_bit_it_3_vnu_108_in_2, msg_to_bit_it_3_vnu_109_in_0, msg_to_bit_it_3_vnu_109_in_1, msg_to_bit_it_3_vnu_109_in_2, msg_to_bit_it_3_vnu_110_in_0, msg_to_bit_it_3_vnu_110_in_1, msg_to_bit_it_3_vnu_110_in_2, msg_to_bit_it_3_vnu_111_in_0, msg_to_bit_it_3_vnu_111_in_1, msg_to_bit_it_3_vnu_111_in_2, msg_to_bit_it_3_vnu_112_in_0, msg_to_bit_it_3_vnu_112_in_1, msg_to_bit_it_3_vnu_112_in_2, msg_to_bit_it_3_vnu_113_in_0, msg_to_bit_it_3_vnu_113_in_1, msg_to_bit_it_3_vnu_113_in_2, msg_to_bit_it_3_vnu_114_in_0, msg_to_bit_it_3_vnu_114_in_1, msg_to_bit_it_3_vnu_114_in_2, msg_to_bit_it_3_vnu_115_in_0, msg_to_bit_it_3_vnu_115_in_1, msg_to_bit_it_3_vnu_115_in_2, msg_to_bit_it_3_vnu_116_in_0, msg_to_bit_it_3_vnu_116_in_1, msg_to_bit_it_3_vnu_116_in_2, msg_to_bit_it_3_vnu_117_in_0, msg_to_bit_it_3_vnu_117_in_1, msg_to_bit_it_3_vnu_117_in_2, msg_to_bit_it_3_vnu_118_in_0, msg_to_bit_it_3_vnu_118_in_1, msg_to_bit_it_3_vnu_118_in_2, msg_to_bit_it_3_vnu_119_in_0, msg_to_bit_it_3_vnu_119_in_1, msg_to_bit_it_3_vnu_119_in_2, msg_to_bit_it_3_vnu_120_in_0, msg_to_bit_it_3_vnu_120_in_1, msg_to_bit_it_3_vnu_120_in_2, msg_to_bit_it_3_vnu_121_in_0, msg_to_bit_it_3_vnu_121_in_1, msg_to_bit_it_3_vnu_121_in_2, msg_to_bit_it_3_vnu_122_in_0, msg_to_bit_it_3_vnu_122_in_1, msg_to_bit_it_3_vnu_122_in_2, msg_to_bit_it_3_vnu_123_in_0, msg_to_bit_it_3_vnu_123_in_1, msg_to_bit_it_3_vnu_123_in_2, msg_to_bit_it_3_vnu_124_in_0, msg_to_bit_it_3_vnu_124_in_1, msg_to_bit_it_3_vnu_124_in_2, msg_to_bit_it_3_vnu_125_in_0, msg_to_bit_it_3_vnu_125_in_1, msg_to_bit_it_3_vnu_125_in_2, msg_to_bit_it_3_vnu_126_in_0, msg_to_bit_it_3_vnu_126_in_1, msg_to_bit_it_3_vnu_126_in_2, msg_to_bit_it_3_vnu_127_in_0, msg_to_bit_it_3_vnu_127_in_1, msg_to_bit_it_3_vnu_127_in_2, msg_to_bit_it_3_vnu_128_in_0, msg_to_bit_it_3_vnu_128_in_1, msg_to_bit_it_3_vnu_128_in_2, msg_to_bit_it_3_vnu_129_in_0, msg_to_bit_it_3_vnu_129_in_1, msg_to_bit_it_3_vnu_129_in_2, msg_to_bit_it_3_vnu_130_in_0, msg_to_bit_it_3_vnu_130_in_1, msg_to_bit_it_3_vnu_130_in_2, msg_to_bit_it_3_vnu_131_in_0, msg_to_bit_it_3_vnu_131_in_1, msg_to_bit_it_3_vnu_131_in_2, msg_to_bit_it_3_vnu_132_in_0, msg_to_bit_it_3_vnu_132_in_1, msg_to_bit_it_3_vnu_132_in_2, msg_to_bit_it_3_vnu_133_in_0, msg_to_bit_it_3_vnu_133_in_1, msg_to_bit_it_3_vnu_133_in_2, msg_to_bit_it_3_vnu_134_in_0, msg_to_bit_it_3_vnu_134_in_1, msg_to_bit_it_3_vnu_134_in_2, msg_to_bit_it_3_vnu_135_in_0, msg_to_bit_it_3_vnu_135_in_1, msg_to_bit_it_3_vnu_135_in_2, msg_to_bit_it_3_vnu_136_in_0, msg_to_bit_it_3_vnu_136_in_1, msg_to_bit_it_3_vnu_136_in_2, msg_to_bit_it_3_vnu_137_in_0, msg_to_bit_it_3_vnu_137_in_1, msg_to_bit_it_3_vnu_137_in_2, msg_to_bit_it_3_vnu_138_in_0, msg_to_bit_it_3_vnu_138_in_1, msg_to_bit_it_3_vnu_138_in_2, msg_to_bit_it_3_vnu_139_in_0, msg_to_bit_it_3_vnu_139_in_1, msg_to_bit_it_3_vnu_139_in_2, msg_to_bit_it_3_vnu_140_in_0, msg_to_bit_it_3_vnu_140_in_1, msg_to_bit_it_3_vnu_140_in_2, msg_to_bit_it_3_vnu_141_in_0, msg_to_bit_it_3_vnu_141_in_1, msg_to_bit_it_3_vnu_141_in_2, msg_to_bit_it_3_vnu_142_in_0, msg_to_bit_it_3_vnu_142_in_1, msg_to_bit_it_3_vnu_142_in_2, msg_to_bit_it_3_vnu_143_in_0, msg_to_bit_it_3_vnu_143_in_1, msg_to_bit_it_3_vnu_143_in_2, msg_to_bit_it_3_vnu_144_in_0, msg_to_bit_it_3_vnu_144_in_1, msg_to_bit_it_3_vnu_144_in_2, msg_to_bit_it_3_vnu_145_in_0, msg_to_bit_it_3_vnu_145_in_1, msg_to_bit_it_3_vnu_145_in_2, msg_to_bit_it_3_vnu_146_in_0, msg_to_bit_it_3_vnu_146_in_1, msg_to_bit_it_3_vnu_146_in_2, msg_to_bit_it_3_vnu_147_in_0, msg_to_bit_it_3_vnu_147_in_1, msg_to_bit_it_3_vnu_147_in_2, msg_to_bit_it_3_vnu_148_in_0, msg_to_bit_it_3_vnu_148_in_1, msg_to_bit_it_3_vnu_148_in_2, msg_to_bit_it_3_vnu_149_in_0, msg_to_bit_it_3_vnu_149_in_1, msg_to_bit_it_3_vnu_149_in_2, msg_to_bit_it_3_vnu_150_in_0, msg_to_bit_it_3_vnu_150_in_1, msg_to_bit_it_3_vnu_150_in_2, msg_to_bit_it_3_vnu_151_in_0, msg_to_bit_it_3_vnu_151_in_1, msg_to_bit_it_3_vnu_151_in_2, msg_to_bit_it_3_vnu_152_in_0, msg_to_bit_it_3_vnu_152_in_1, msg_to_bit_it_3_vnu_152_in_2, msg_to_bit_it_3_vnu_153_in_0, msg_to_bit_it_3_vnu_153_in_1, msg_to_bit_it_3_vnu_153_in_2, msg_to_bit_it_3_vnu_154_in_0, msg_to_bit_it_3_vnu_154_in_1, msg_to_bit_it_3_vnu_154_in_2, msg_to_bit_it_3_vnu_155_in_0, msg_to_bit_it_3_vnu_155_in_1, msg_to_bit_it_3_vnu_155_in_2, msg_to_bit_it_3_vnu_156_in_0, msg_to_bit_it_3_vnu_156_in_1, msg_to_bit_it_3_vnu_156_in_2, msg_to_bit_it_3_vnu_157_in_0, msg_to_bit_it_3_vnu_157_in_1, msg_to_bit_it_3_vnu_157_in_2, msg_to_bit_it_3_vnu_158_in_0, msg_to_bit_it_3_vnu_158_in_1, msg_to_bit_it_3_vnu_158_in_2, msg_to_bit_it_3_vnu_159_in_0, msg_to_bit_it_3_vnu_159_in_1, msg_to_bit_it_3_vnu_159_in_2, msg_to_bit_it_3_vnu_160_in_0, msg_to_bit_it_3_vnu_160_in_1, msg_to_bit_it_3_vnu_160_in_2, msg_to_bit_it_3_vnu_161_in_0, msg_to_bit_it_3_vnu_161_in_1, msg_to_bit_it_3_vnu_161_in_2, msg_to_bit_it_3_vnu_162_in_0, msg_to_bit_it_3_vnu_162_in_1, msg_to_bit_it_3_vnu_162_in_2, msg_to_bit_it_3_vnu_163_in_0, msg_to_bit_it_3_vnu_163_in_1, msg_to_bit_it_3_vnu_163_in_2, msg_to_bit_it_3_vnu_164_in_0, msg_to_bit_it_3_vnu_164_in_1, msg_to_bit_it_3_vnu_164_in_2, msg_to_bit_it_3_vnu_165_in_0, msg_to_bit_it_3_vnu_165_in_1, msg_to_bit_it_3_vnu_165_in_2, msg_to_bit_it_3_vnu_166_in_0, msg_to_bit_it_3_vnu_166_in_1, msg_to_bit_it_3_vnu_166_in_2, msg_to_bit_it_3_vnu_167_in_0, msg_to_bit_it_3_vnu_167_in_1, msg_to_bit_it_3_vnu_167_in_2, msg_to_bit_it_3_vnu_168_in_0, msg_to_bit_it_3_vnu_168_in_1, msg_to_bit_it_3_vnu_168_in_2, msg_to_bit_it_3_vnu_169_in_0, msg_to_bit_it_3_vnu_169_in_1, msg_to_bit_it_3_vnu_169_in_2, msg_to_bit_it_3_vnu_170_in_0, msg_to_bit_it_3_vnu_170_in_1, msg_to_bit_it_3_vnu_170_in_2, msg_to_bit_it_3_vnu_171_in_0, msg_to_bit_it_3_vnu_171_in_1, msg_to_bit_it_3_vnu_171_in_2, msg_to_bit_it_3_vnu_172_in_0, msg_to_bit_it_3_vnu_172_in_1, msg_to_bit_it_3_vnu_172_in_2, msg_to_bit_it_3_vnu_173_in_0, msg_to_bit_it_3_vnu_173_in_1, msg_to_bit_it_3_vnu_173_in_2, msg_to_bit_it_3_vnu_174_in_0, msg_to_bit_it_3_vnu_174_in_1, msg_to_bit_it_3_vnu_174_in_2, msg_to_bit_it_3_vnu_175_in_0, msg_to_bit_it_3_vnu_175_in_1, msg_to_bit_it_3_vnu_175_in_2, msg_to_bit_it_3_vnu_176_in_0, msg_to_bit_it_3_vnu_176_in_1, msg_to_bit_it_3_vnu_176_in_2, msg_to_bit_it_3_vnu_177_in_0, msg_to_bit_it_3_vnu_177_in_1, msg_to_bit_it_3_vnu_177_in_2, msg_to_bit_it_3_vnu_178_in_0, msg_to_bit_it_3_vnu_178_in_1, msg_to_bit_it_3_vnu_178_in_2, msg_to_bit_it_3_vnu_179_in_0, msg_to_bit_it_3_vnu_179_in_1, msg_to_bit_it_3_vnu_179_in_2, msg_to_bit_it_3_vnu_180_in_0, msg_to_bit_it_3_vnu_180_in_1, msg_to_bit_it_3_vnu_180_in_2, msg_to_bit_it_3_vnu_181_in_0, msg_to_bit_it_3_vnu_181_in_1, msg_to_bit_it_3_vnu_181_in_2, msg_to_bit_it_3_vnu_182_in_0, msg_to_bit_it_3_vnu_182_in_1, msg_to_bit_it_3_vnu_182_in_2, msg_to_bit_it_3_vnu_183_in_0, msg_to_bit_it_3_vnu_183_in_1, msg_to_bit_it_3_vnu_183_in_2, msg_to_bit_it_3_vnu_184_in_0, msg_to_bit_it_3_vnu_184_in_1, msg_to_bit_it_3_vnu_184_in_2, msg_to_bit_it_3_vnu_185_in_0, msg_to_bit_it_3_vnu_185_in_1, msg_to_bit_it_3_vnu_185_in_2, msg_to_bit_it_3_vnu_186_in_0, msg_to_bit_it_3_vnu_186_in_1, msg_to_bit_it_3_vnu_186_in_2, msg_to_bit_it_3_vnu_187_in_0, msg_to_bit_it_3_vnu_187_in_1, msg_to_bit_it_3_vnu_187_in_2, msg_to_bit_it_3_vnu_188_in_0, msg_to_bit_it_3_vnu_188_in_1, msg_to_bit_it_3_vnu_188_in_2, msg_to_bit_it_3_vnu_189_in_0, msg_to_bit_it_3_vnu_189_in_1, msg_to_bit_it_3_vnu_189_in_2, msg_to_bit_it_3_vnu_190_in_0, msg_to_bit_it_3_vnu_190_in_1, msg_to_bit_it_3_vnu_190_in_2, msg_to_bit_it_3_vnu_191_in_0, msg_to_bit_it_3_vnu_191_in_1, msg_to_bit_it_3_vnu_191_in_2, msg_to_bit_it_3_vnu_192_in_0, msg_to_bit_it_3_vnu_192_in_1, msg_to_bit_it_3_vnu_192_in_2, msg_to_bit_it_3_vnu_193_in_0, msg_to_bit_it_3_vnu_193_in_1, msg_to_bit_it_3_vnu_193_in_2, msg_to_bit_it_3_vnu_194_in_0, msg_to_bit_it_3_vnu_194_in_1, msg_to_bit_it_3_vnu_194_in_2, msg_to_bit_it_3_vnu_195_in_0, msg_to_bit_it_3_vnu_195_in_1, msg_to_bit_it_3_vnu_195_in_2, msg_to_bit_it_3_vnu_196_in_0, msg_to_bit_it_3_vnu_196_in_1, msg_to_bit_it_3_vnu_196_in_2, msg_to_bit_it_3_vnu_197_in_0, msg_to_bit_it_3_vnu_197_in_1, msg_to_bit_it_3_vnu_197_in_2, msg_to_bit_it_4_vnu_0_in_0, msg_to_bit_it_4_vnu_0_in_1, msg_to_bit_it_4_vnu_0_in_2, msg_to_bit_it_4_vnu_1_in_0, msg_to_bit_it_4_vnu_1_in_1, msg_to_bit_it_4_vnu_1_in_2, msg_to_bit_it_4_vnu_2_in_0, msg_to_bit_it_4_vnu_2_in_1, msg_to_bit_it_4_vnu_2_in_2, msg_to_bit_it_4_vnu_3_in_0, msg_to_bit_it_4_vnu_3_in_1, msg_to_bit_it_4_vnu_3_in_2, msg_to_bit_it_4_vnu_4_in_0, msg_to_bit_it_4_vnu_4_in_1, msg_to_bit_it_4_vnu_4_in_2, msg_to_bit_it_4_vnu_5_in_0, msg_to_bit_it_4_vnu_5_in_1, msg_to_bit_it_4_vnu_5_in_2, msg_to_bit_it_4_vnu_6_in_0, msg_to_bit_it_4_vnu_6_in_1, msg_to_bit_it_4_vnu_6_in_2, msg_to_bit_it_4_vnu_7_in_0, msg_to_bit_it_4_vnu_7_in_1, msg_to_bit_it_4_vnu_7_in_2, msg_to_bit_it_4_vnu_8_in_0, msg_to_bit_it_4_vnu_8_in_1, msg_to_bit_it_4_vnu_8_in_2, msg_to_bit_it_4_vnu_9_in_0, msg_to_bit_it_4_vnu_9_in_1, msg_to_bit_it_4_vnu_9_in_2, msg_to_bit_it_4_vnu_10_in_0, msg_to_bit_it_4_vnu_10_in_1, msg_to_bit_it_4_vnu_10_in_2, msg_to_bit_it_4_vnu_11_in_0, msg_to_bit_it_4_vnu_11_in_1, msg_to_bit_it_4_vnu_11_in_2, msg_to_bit_it_4_vnu_12_in_0, msg_to_bit_it_4_vnu_12_in_1, msg_to_bit_it_4_vnu_12_in_2, msg_to_bit_it_4_vnu_13_in_0, msg_to_bit_it_4_vnu_13_in_1, msg_to_bit_it_4_vnu_13_in_2, msg_to_bit_it_4_vnu_14_in_0, msg_to_bit_it_4_vnu_14_in_1, msg_to_bit_it_4_vnu_14_in_2, msg_to_bit_it_4_vnu_15_in_0, msg_to_bit_it_4_vnu_15_in_1, msg_to_bit_it_4_vnu_15_in_2, msg_to_bit_it_4_vnu_16_in_0, msg_to_bit_it_4_vnu_16_in_1, msg_to_bit_it_4_vnu_16_in_2, msg_to_bit_it_4_vnu_17_in_0, msg_to_bit_it_4_vnu_17_in_1, msg_to_bit_it_4_vnu_17_in_2, msg_to_bit_it_4_vnu_18_in_0, msg_to_bit_it_4_vnu_18_in_1, msg_to_bit_it_4_vnu_18_in_2, msg_to_bit_it_4_vnu_19_in_0, msg_to_bit_it_4_vnu_19_in_1, msg_to_bit_it_4_vnu_19_in_2, msg_to_bit_it_4_vnu_20_in_0, msg_to_bit_it_4_vnu_20_in_1, msg_to_bit_it_4_vnu_20_in_2, msg_to_bit_it_4_vnu_21_in_0, msg_to_bit_it_4_vnu_21_in_1, msg_to_bit_it_4_vnu_21_in_2, msg_to_bit_it_4_vnu_22_in_0, msg_to_bit_it_4_vnu_22_in_1, msg_to_bit_it_4_vnu_22_in_2, msg_to_bit_it_4_vnu_23_in_0, msg_to_bit_it_4_vnu_23_in_1, msg_to_bit_it_4_vnu_23_in_2, msg_to_bit_it_4_vnu_24_in_0, msg_to_bit_it_4_vnu_24_in_1, msg_to_bit_it_4_vnu_24_in_2, msg_to_bit_it_4_vnu_25_in_0, msg_to_bit_it_4_vnu_25_in_1, msg_to_bit_it_4_vnu_25_in_2, msg_to_bit_it_4_vnu_26_in_0, msg_to_bit_it_4_vnu_26_in_1, msg_to_bit_it_4_vnu_26_in_2, msg_to_bit_it_4_vnu_27_in_0, msg_to_bit_it_4_vnu_27_in_1, msg_to_bit_it_4_vnu_27_in_2, msg_to_bit_it_4_vnu_28_in_0, msg_to_bit_it_4_vnu_28_in_1, msg_to_bit_it_4_vnu_28_in_2, msg_to_bit_it_4_vnu_29_in_0, msg_to_bit_it_4_vnu_29_in_1, msg_to_bit_it_4_vnu_29_in_2, msg_to_bit_it_4_vnu_30_in_0, msg_to_bit_it_4_vnu_30_in_1, msg_to_bit_it_4_vnu_30_in_2, msg_to_bit_it_4_vnu_31_in_0, msg_to_bit_it_4_vnu_31_in_1, msg_to_bit_it_4_vnu_31_in_2, msg_to_bit_it_4_vnu_32_in_0, msg_to_bit_it_4_vnu_32_in_1, msg_to_bit_it_4_vnu_32_in_2, msg_to_bit_it_4_vnu_33_in_0, msg_to_bit_it_4_vnu_33_in_1, msg_to_bit_it_4_vnu_33_in_2, msg_to_bit_it_4_vnu_34_in_0, msg_to_bit_it_4_vnu_34_in_1, msg_to_bit_it_4_vnu_34_in_2, msg_to_bit_it_4_vnu_35_in_0, msg_to_bit_it_4_vnu_35_in_1, msg_to_bit_it_4_vnu_35_in_2, msg_to_bit_it_4_vnu_36_in_0, msg_to_bit_it_4_vnu_36_in_1, msg_to_bit_it_4_vnu_36_in_2, msg_to_bit_it_4_vnu_37_in_0, msg_to_bit_it_4_vnu_37_in_1, msg_to_bit_it_4_vnu_37_in_2, msg_to_bit_it_4_vnu_38_in_0, msg_to_bit_it_4_vnu_38_in_1, msg_to_bit_it_4_vnu_38_in_2, msg_to_bit_it_4_vnu_39_in_0, msg_to_bit_it_4_vnu_39_in_1, msg_to_bit_it_4_vnu_39_in_2, msg_to_bit_it_4_vnu_40_in_0, msg_to_bit_it_4_vnu_40_in_1, msg_to_bit_it_4_vnu_40_in_2, msg_to_bit_it_4_vnu_41_in_0, msg_to_bit_it_4_vnu_41_in_1, msg_to_bit_it_4_vnu_41_in_2, msg_to_bit_it_4_vnu_42_in_0, msg_to_bit_it_4_vnu_42_in_1, msg_to_bit_it_4_vnu_42_in_2, msg_to_bit_it_4_vnu_43_in_0, msg_to_bit_it_4_vnu_43_in_1, msg_to_bit_it_4_vnu_43_in_2, msg_to_bit_it_4_vnu_44_in_0, msg_to_bit_it_4_vnu_44_in_1, msg_to_bit_it_4_vnu_44_in_2, msg_to_bit_it_4_vnu_45_in_0, msg_to_bit_it_4_vnu_45_in_1, msg_to_bit_it_4_vnu_45_in_2, msg_to_bit_it_4_vnu_46_in_0, msg_to_bit_it_4_vnu_46_in_1, msg_to_bit_it_4_vnu_46_in_2, msg_to_bit_it_4_vnu_47_in_0, msg_to_bit_it_4_vnu_47_in_1, msg_to_bit_it_4_vnu_47_in_2, msg_to_bit_it_4_vnu_48_in_0, msg_to_bit_it_4_vnu_48_in_1, msg_to_bit_it_4_vnu_48_in_2, msg_to_bit_it_4_vnu_49_in_0, msg_to_bit_it_4_vnu_49_in_1, msg_to_bit_it_4_vnu_49_in_2, msg_to_bit_it_4_vnu_50_in_0, msg_to_bit_it_4_vnu_50_in_1, msg_to_bit_it_4_vnu_50_in_2, msg_to_bit_it_4_vnu_51_in_0, msg_to_bit_it_4_vnu_51_in_1, msg_to_bit_it_4_vnu_51_in_2, msg_to_bit_it_4_vnu_52_in_0, msg_to_bit_it_4_vnu_52_in_1, msg_to_bit_it_4_vnu_52_in_2, msg_to_bit_it_4_vnu_53_in_0, msg_to_bit_it_4_vnu_53_in_1, msg_to_bit_it_4_vnu_53_in_2, msg_to_bit_it_4_vnu_54_in_0, msg_to_bit_it_4_vnu_54_in_1, msg_to_bit_it_4_vnu_54_in_2, msg_to_bit_it_4_vnu_55_in_0, msg_to_bit_it_4_vnu_55_in_1, msg_to_bit_it_4_vnu_55_in_2, msg_to_bit_it_4_vnu_56_in_0, msg_to_bit_it_4_vnu_56_in_1, msg_to_bit_it_4_vnu_56_in_2, msg_to_bit_it_4_vnu_57_in_0, msg_to_bit_it_4_vnu_57_in_1, msg_to_bit_it_4_vnu_57_in_2, msg_to_bit_it_4_vnu_58_in_0, msg_to_bit_it_4_vnu_58_in_1, msg_to_bit_it_4_vnu_58_in_2, msg_to_bit_it_4_vnu_59_in_0, msg_to_bit_it_4_vnu_59_in_1, msg_to_bit_it_4_vnu_59_in_2, msg_to_bit_it_4_vnu_60_in_0, msg_to_bit_it_4_vnu_60_in_1, msg_to_bit_it_4_vnu_60_in_2, msg_to_bit_it_4_vnu_61_in_0, msg_to_bit_it_4_vnu_61_in_1, msg_to_bit_it_4_vnu_61_in_2, msg_to_bit_it_4_vnu_62_in_0, msg_to_bit_it_4_vnu_62_in_1, msg_to_bit_it_4_vnu_62_in_2, msg_to_bit_it_4_vnu_63_in_0, msg_to_bit_it_4_vnu_63_in_1, msg_to_bit_it_4_vnu_63_in_2, msg_to_bit_it_4_vnu_64_in_0, msg_to_bit_it_4_vnu_64_in_1, msg_to_bit_it_4_vnu_64_in_2, msg_to_bit_it_4_vnu_65_in_0, msg_to_bit_it_4_vnu_65_in_1, msg_to_bit_it_4_vnu_65_in_2, msg_to_bit_it_4_vnu_66_in_0, msg_to_bit_it_4_vnu_66_in_1, msg_to_bit_it_4_vnu_66_in_2, msg_to_bit_it_4_vnu_67_in_0, msg_to_bit_it_4_vnu_67_in_1, msg_to_bit_it_4_vnu_67_in_2, msg_to_bit_it_4_vnu_68_in_0, msg_to_bit_it_4_vnu_68_in_1, msg_to_bit_it_4_vnu_68_in_2, msg_to_bit_it_4_vnu_69_in_0, msg_to_bit_it_4_vnu_69_in_1, msg_to_bit_it_4_vnu_69_in_2, msg_to_bit_it_4_vnu_70_in_0, msg_to_bit_it_4_vnu_70_in_1, msg_to_bit_it_4_vnu_70_in_2, msg_to_bit_it_4_vnu_71_in_0, msg_to_bit_it_4_vnu_71_in_1, msg_to_bit_it_4_vnu_71_in_2, msg_to_bit_it_4_vnu_72_in_0, msg_to_bit_it_4_vnu_72_in_1, msg_to_bit_it_4_vnu_72_in_2, msg_to_bit_it_4_vnu_73_in_0, msg_to_bit_it_4_vnu_73_in_1, msg_to_bit_it_4_vnu_73_in_2, msg_to_bit_it_4_vnu_74_in_0, msg_to_bit_it_4_vnu_74_in_1, msg_to_bit_it_4_vnu_74_in_2, msg_to_bit_it_4_vnu_75_in_0, msg_to_bit_it_4_vnu_75_in_1, msg_to_bit_it_4_vnu_75_in_2, msg_to_bit_it_4_vnu_76_in_0, msg_to_bit_it_4_vnu_76_in_1, msg_to_bit_it_4_vnu_76_in_2, msg_to_bit_it_4_vnu_77_in_0, msg_to_bit_it_4_vnu_77_in_1, msg_to_bit_it_4_vnu_77_in_2, msg_to_bit_it_4_vnu_78_in_0, msg_to_bit_it_4_vnu_78_in_1, msg_to_bit_it_4_vnu_78_in_2, msg_to_bit_it_4_vnu_79_in_0, msg_to_bit_it_4_vnu_79_in_1, msg_to_bit_it_4_vnu_79_in_2, msg_to_bit_it_4_vnu_80_in_0, msg_to_bit_it_4_vnu_80_in_1, msg_to_bit_it_4_vnu_80_in_2, msg_to_bit_it_4_vnu_81_in_0, msg_to_bit_it_4_vnu_81_in_1, msg_to_bit_it_4_vnu_81_in_2, msg_to_bit_it_4_vnu_82_in_0, msg_to_bit_it_4_vnu_82_in_1, msg_to_bit_it_4_vnu_82_in_2, msg_to_bit_it_4_vnu_83_in_0, msg_to_bit_it_4_vnu_83_in_1, msg_to_bit_it_4_vnu_83_in_2, msg_to_bit_it_4_vnu_84_in_0, msg_to_bit_it_4_vnu_84_in_1, msg_to_bit_it_4_vnu_84_in_2, msg_to_bit_it_4_vnu_85_in_0, msg_to_bit_it_4_vnu_85_in_1, msg_to_bit_it_4_vnu_85_in_2, msg_to_bit_it_4_vnu_86_in_0, msg_to_bit_it_4_vnu_86_in_1, msg_to_bit_it_4_vnu_86_in_2, msg_to_bit_it_4_vnu_87_in_0, msg_to_bit_it_4_vnu_87_in_1, msg_to_bit_it_4_vnu_87_in_2, msg_to_bit_it_4_vnu_88_in_0, msg_to_bit_it_4_vnu_88_in_1, msg_to_bit_it_4_vnu_88_in_2, msg_to_bit_it_4_vnu_89_in_0, msg_to_bit_it_4_vnu_89_in_1, msg_to_bit_it_4_vnu_89_in_2, msg_to_bit_it_4_vnu_90_in_0, msg_to_bit_it_4_vnu_90_in_1, msg_to_bit_it_4_vnu_90_in_2, msg_to_bit_it_4_vnu_91_in_0, msg_to_bit_it_4_vnu_91_in_1, msg_to_bit_it_4_vnu_91_in_2, msg_to_bit_it_4_vnu_92_in_0, msg_to_bit_it_4_vnu_92_in_1, msg_to_bit_it_4_vnu_92_in_2, msg_to_bit_it_4_vnu_93_in_0, msg_to_bit_it_4_vnu_93_in_1, msg_to_bit_it_4_vnu_93_in_2, msg_to_bit_it_4_vnu_94_in_0, msg_to_bit_it_4_vnu_94_in_1, msg_to_bit_it_4_vnu_94_in_2, msg_to_bit_it_4_vnu_95_in_0, msg_to_bit_it_4_vnu_95_in_1, msg_to_bit_it_4_vnu_95_in_2, msg_to_bit_it_4_vnu_96_in_0, msg_to_bit_it_4_vnu_96_in_1, msg_to_bit_it_4_vnu_96_in_2, msg_to_bit_it_4_vnu_97_in_0, msg_to_bit_it_4_vnu_97_in_1, msg_to_bit_it_4_vnu_97_in_2, msg_to_bit_it_4_vnu_98_in_0, msg_to_bit_it_4_vnu_98_in_1, msg_to_bit_it_4_vnu_98_in_2, msg_to_bit_it_4_vnu_99_in_0, msg_to_bit_it_4_vnu_99_in_1, msg_to_bit_it_4_vnu_99_in_2, msg_to_bit_it_4_vnu_100_in_0, msg_to_bit_it_4_vnu_100_in_1, msg_to_bit_it_4_vnu_100_in_2, msg_to_bit_it_4_vnu_101_in_0, msg_to_bit_it_4_vnu_101_in_1, msg_to_bit_it_4_vnu_101_in_2, msg_to_bit_it_4_vnu_102_in_0, msg_to_bit_it_4_vnu_102_in_1, msg_to_bit_it_4_vnu_102_in_2, msg_to_bit_it_4_vnu_103_in_0, msg_to_bit_it_4_vnu_103_in_1, msg_to_bit_it_4_vnu_103_in_2, msg_to_bit_it_4_vnu_104_in_0, msg_to_bit_it_4_vnu_104_in_1, msg_to_bit_it_4_vnu_104_in_2, msg_to_bit_it_4_vnu_105_in_0, msg_to_bit_it_4_vnu_105_in_1, msg_to_bit_it_4_vnu_105_in_2, msg_to_bit_it_4_vnu_106_in_0, msg_to_bit_it_4_vnu_106_in_1, msg_to_bit_it_4_vnu_106_in_2, msg_to_bit_it_4_vnu_107_in_0, msg_to_bit_it_4_vnu_107_in_1, msg_to_bit_it_4_vnu_107_in_2, msg_to_bit_it_4_vnu_108_in_0, msg_to_bit_it_4_vnu_108_in_1, msg_to_bit_it_4_vnu_108_in_2, msg_to_bit_it_4_vnu_109_in_0, msg_to_bit_it_4_vnu_109_in_1, msg_to_bit_it_4_vnu_109_in_2, msg_to_bit_it_4_vnu_110_in_0, msg_to_bit_it_4_vnu_110_in_1, msg_to_bit_it_4_vnu_110_in_2, msg_to_bit_it_4_vnu_111_in_0, msg_to_bit_it_4_vnu_111_in_1, msg_to_bit_it_4_vnu_111_in_2, msg_to_bit_it_4_vnu_112_in_0, msg_to_bit_it_4_vnu_112_in_1, msg_to_bit_it_4_vnu_112_in_2, msg_to_bit_it_4_vnu_113_in_0, msg_to_bit_it_4_vnu_113_in_1, msg_to_bit_it_4_vnu_113_in_2, msg_to_bit_it_4_vnu_114_in_0, msg_to_bit_it_4_vnu_114_in_1, msg_to_bit_it_4_vnu_114_in_2, msg_to_bit_it_4_vnu_115_in_0, msg_to_bit_it_4_vnu_115_in_1, msg_to_bit_it_4_vnu_115_in_2, msg_to_bit_it_4_vnu_116_in_0, msg_to_bit_it_4_vnu_116_in_1, msg_to_bit_it_4_vnu_116_in_2, msg_to_bit_it_4_vnu_117_in_0, msg_to_bit_it_4_vnu_117_in_1, msg_to_bit_it_4_vnu_117_in_2, msg_to_bit_it_4_vnu_118_in_0, msg_to_bit_it_4_vnu_118_in_1, msg_to_bit_it_4_vnu_118_in_2, msg_to_bit_it_4_vnu_119_in_0, msg_to_bit_it_4_vnu_119_in_1, msg_to_bit_it_4_vnu_119_in_2, msg_to_bit_it_4_vnu_120_in_0, msg_to_bit_it_4_vnu_120_in_1, msg_to_bit_it_4_vnu_120_in_2, msg_to_bit_it_4_vnu_121_in_0, msg_to_bit_it_4_vnu_121_in_1, msg_to_bit_it_4_vnu_121_in_2, msg_to_bit_it_4_vnu_122_in_0, msg_to_bit_it_4_vnu_122_in_1, msg_to_bit_it_4_vnu_122_in_2, msg_to_bit_it_4_vnu_123_in_0, msg_to_bit_it_4_vnu_123_in_1, msg_to_bit_it_4_vnu_123_in_2, msg_to_bit_it_4_vnu_124_in_0, msg_to_bit_it_4_vnu_124_in_1, msg_to_bit_it_4_vnu_124_in_2, msg_to_bit_it_4_vnu_125_in_0, msg_to_bit_it_4_vnu_125_in_1, msg_to_bit_it_4_vnu_125_in_2, msg_to_bit_it_4_vnu_126_in_0, msg_to_bit_it_4_vnu_126_in_1, msg_to_bit_it_4_vnu_126_in_2, msg_to_bit_it_4_vnu_127_in_0, msg_to_bit_it_4_vnu_127_in_1, msg_to_bit_it_4_vnu_127_in_2, msg_to_bit_it_4_vnu_128_in_0, msg_to_bit_it_4_vnu_128_in_1, msg_to_bit_it_4_vnu_128_in_2, msg_to_bit_it_4_vnu_129_in_0, msg_to_bit_it_4_vnu_129_in_1, msg_to_bit_it_4_vnu_129_in_2, msg_to_bit_it_4_vnu_130_in_0, msg_to_bit_it_4_vnu_130_in_1, msg_to_bit_it_4_vnu_130_in_2, msg_to_bit_it_4_vnu_131_in_0, msg_to_bit_it_4_vnu_131_in_1, msg_to_bit_it_4_vnu_131_in_2, msg_to_bit_it_4_vnu_132_in_0, msg_to_bit_it_4_vnu_132_in_1, msg_to_bit_it_4_vnu_132_in_2, msg_to_bit_it_4_vnu_133_in_0, msg_to_bit_it_4_vnu_133_in_1, msg_to_bit_it_4_vnu_133_in_2, msg_to_bit_it_4_vnu_134_in_0, msg_to_bit_it_4_vnu_134_in_1, msg_to_bit_it_4_vnu_134_in_2, msg_to_bit_it_4_vnu_135_in_0, msg_to_bit_it_4_vnu_135_in_1, msg_to_bit_it_4_vnu_135_in_2, msg_to_bit_it_4_vnu_136_in_0, msg_to_bit_it_4_vnu_136_in_1, msg_to_bit_it_4_vnu_136_in_2, msg_to_bit_it_4_vnu_137_in_0, msg_to_bit_it_4_vnu_137_in_1, msg_to_bit_it_4_vnu_137_in_2, msg_to_bit_it_4_vnu_138_in_0, msg_to_bit_it_4_vnu_138_in_1, msg_to_bit_it_4_vnu_138_in_2, msg_to_bit_it_4_vnu_139_in_0, msg_to_bit_it_4_vnu_139_in_1, msg_to_bit_it_4_vnu_139_in_2, msg_to_bit_it_4_vnu_140_in_0, msg_to_bit_it_4_vnu_140_in_1, msg_to_bit_it_4_vnu_140_in_2, msg_to_bit_it_4_vnu_141_in_0, msg_to_bit_it_4_vnu_141_in_1, msg_to_bit_it_4_vnu_141_in_2, msg_to_bit_it_4_vnu_142_in_0, msg_to_bit_it_4_vnu_142_in_1, msg_to_bit_it_4_vnu_142_in_2, msg_to_bit_it_4_vnu_143_in_0, msg_to_bit_it_4_vnu_143_in_1, msg_to_bit_it_4_vnu_143_in_2, msg_to_bit_it_4_vnu_144_in_0, msg_to_bit_it_4_vnu_144_in_1, msg_to_bit_it_4_vnu_144_in_2, msg_to_bit_it_4_vnu_145_in_0, msg_to_bit_it_4_vnu_145_in_1, msg_to_bit_it_4_vnu_145_in_2, msg_to_bit_it_4_vnu_146_in_0, msg_to_bit_it_4_vnu_146_in_1, msg_to_bit_it_4_vnu_146_in_2, msg_to_bit_it_4_vnu_147_in_0, msg_to_bit_it_4_vnu_147_in_1, msg_to_bit_it_4_vnu_147_in_2, msg_to_bit_it_4_vnu_148_in_0, msg_to_bit_it_4_vnu_148_in_1, msg_to_bit_it_4_vnu_148_in_2, msg_to_bit_it_4_vnu_149_in_0, msg_to_bit_it_4_vnu_149_in_1, msg_to_bit_it_4_vnu_149_in_2, msg_to_bit_it_4_vnu_150_in_0, msg_to_bit_it_4_vnu_150_in_1, msg_to_bit_it_4_vnu_150_in_2, msg_to_bit_it_4_vnu_151_in_0, msg_to_bit_it_4_vnu_151_in_1, msg_to_bit_it_4_vnu_151_in_2, msg_to_bit_it_4_vnu_152_in_0, msg_to_bit_it_4_vnu_152_in_1, msg_to_bit_it_4_vnu_152_in_2, msg_to_bit_it_4_vnu_153_in_0, msg_to_bit_it_4_vnu_153_in_1, msg_to_bit_it_4_vnu_153_in_2, msg_to_bit_it_4_vnu_154_in_0, msg_to_bit_it_4_vnu_154_in_1, msg_to_bit_it_4_vnu_154_in_2, msg_to_bit_it_4_vnu_155_in_0, msg_to_bit_it_4_vnu_155_in_1, msg_to_bit_it_4_vnu_155_in_2, msg_to_bit_it_4_vnu_156_in_0, msg_to_bit_it_4_vnu_156_in_1, msg_to_bit_it_4_vnu_156_in_2, msg_to_bit_it_4_vnu_157_in_0, msg_to_bit_it_4_vnu_157_in_1, msg_to_bit_it_4_vnu_157_in_2, msg_to_bit_it_4_vnu_158_in_0, msg_to_bit_it_4_vnu_158_in_1, msg_to_bit_it_4_vnu_158_in_2, msg_to_bit_it_4_vnu_159_in_0, msg_to_bit_it_4_vnu_159_in_1, msg_to_bit_it_4_vnu_159_in_2, msg_to_bit_it_4_vnu_160_in_0, msg_to_bit_it_4_vnu_160_in_1, msg_to_bit_it_4_vnu_160_in_2, msg_to_bit_it_4_vnu_161_in_0, msg_to_bit_it_4_vnu_161_in_1, msg_to_bit_it_4_vnu_161_in_2, msg_to_bit_it_4_vnu_162_in_0, msg_to_bit_it_4_vnu_162_in_1, msg_to_bit_it_4_vnu_162_in_2, msg_to_bit_it_4_vnu_163_in_0, msg_to_bit_it_4_vnu_163_in_1, msg_to_bit_it_4_vnu_163_in_2, msg_to_bit_it_4_vnu_164_in_0, msg_to_bit_it_4_vnu_164_in_1, msg_to_bit_it_4_vnu_164_in_2, msg_to_bit_it_4_vnu_165_in_0, msg_to_bit_it_4_vnu_165_in_1, msg_to_bit_it_4_vnu_165_in_2, msg_to_bit_it_4_vnu_166_in_0, msg_to_bit_it_4_vnu_166_in_1, msg_to_bit_it_4_vnu_166_in_2, msg_to_bit_it_4_vnu_167_in_0, msg_to_bit_it_4_vnu_167_in_1, msg_to_bit_it_4_vnu_167_in_2, msg_to_bit_it_4_vnu_168_in_0, msg_to_bit_it_4_vnu_168_in_1, msg_to_bit_it_4_vnu_168_in_2, msg_to_bit_it_4_vnu_169_in_0, msg_to_bit_it_4_vnu_169_in_1, msg_to_bit_it_4_vnu_169_in_2, msg_to_bit_it_4_vnu_170_in_0, msg_to_bit_it_4_vnu_170_in_1, msg_to_bit_it_4_vnu_170_in_2, msg_to_bit_it_4_vnu_171_in_0, msg_to_bit_it_4_vnu_171_in_1, msg_to_bit_it_4_vnu_171_in_2, msg_to_bit_it_4_vnu_172_in_0, msg_to_bit_it_4_vnu_172_in_1, msg_to_bit_it_4_vnu_172_in_2, msg_to_bit_it_4_vnu_173_in_0, msg_to_bit_it_4_vnu_173_in_1, msg_to_bit_it_4_vnu_173_in_2, msg_to_bit_it_4_vnu_174_in_0, msg_to_bit_it_4_vnu_174_in_1, msg_to_bit_it_4_vnu_174_in_2, msg_to_bit_it_4_vnu_175_in_0, msg_to_bit_it_4_vnu_175_in_1, msg_to_bit_it_4_vnu_175_in_2, msg_to_bit_it_4_vnu_176_in_0, msg_to_bit_it_4_vnu_176_in_1, msg_to_bit_it_4_vnu_176_in_2, msg_to_bit_it_4_vnu_177_in_0, msg_to_bit_it_4_vnu_177_in_1, msg_to_bit_it_4_vnu_177_in_2, msg_to_bit_it_4_vnu_178_in_0, msg_to_bit_it_4_vnu_178_in_1, msg_to_bit_it_4_vnu_178_in_2, msg_to_bit_it_4_vnu_179_in_0, msg_to_bit_it_4_vnu_179_in_1, msg_to_bit_it_4_vnu_179_in_2, msg_to_bit_it_4_vnu_180_in_0, msg_to_bit_it_4_vnu_180_in_1, msg_to_bit_it_4_vnu_180_in_2, msg_to_bit_it_4_vnu_181_in_0, msg_to_bit_it_4_vnu_181_in_1, msg_to_bit_it_4_vnu_181_in_2, msg_to_bit_it_4_vnu_182_in_0, msg_to_bit_it_4_vnu_182_in_1, msg_to_bit_it_4_vnu_182_in_2, msg_to_bit_it_4_vnu_183_in_0, msg_to_bit_it_4_vnu_183_in_1, msg_to_bit_it_4_vnu_183_in_2, msg_to_bit_it_4_vnu_184_in_0, msg_to_bit_it_4_vnu_184_in_1, msg_to_bit_it_4_vnu_184_in_2, msg_to_bit_it_4_vnu_185_in_0, msg_to_bit_it_4_vnu_185_in_1, msg_to_bit_it_4_vnu_185_in_2, msg_to_bit_it_4_vnu_186_in_0, msg_to_bit_it_4_vnu_186_in_1, msg_to_bit_it_4_vnu_186_in_2, msg_to_bit_it_4_vnu_187_in_0, msg_to_bit_it_4_vnu_187_in_1, msg_to_bit_it_4_vnu_187_in_2, msg_to_bit_it_4_vnu_188_in_0, msg_to_bit_it_4_vnu_188_in_1, msg_to_bit_it_4_vnu_188_in_2, msg_to_bit_it_4_vnu_189_in_0, msg_to_bit_it_4_vnu_189_in_1, msg_to_bit_it_4_vnu_189_in_2, msg_to_bit_it_4_vnu_190_in_0, msg_to_bit_it_4_vnu_190_in_1, msg_to_bit_it_4_vnu_190_in_2, msg_to_bit_it_4_vnu_191_in_0, msg_to_bit_it_4_vnu_191_in_1, msg_to_bit_it_4_vnu_191_in_2, msg_to_bit_it_4_vnu_192_in_0, msg_to_bit_it_4_vnu_192_in_1, msg_to_bit_it_4_vnu_192_in_2, msg_to_bit_it_4_vnu_193_in_0, msg_to_bit_it_4_vnu_193_in_1, msg_to_bit_it_4_vnu_193_in_2, msg_to_bit_it_4_vnu_194_in_0, msg_to_bit_it_4_vnu_194_in_1, msg_to_bit_it_4_vnu_194_in_2, msg_to_bit_it_4_vnu_195_in_0, msg_to_bit_it_4_vnu_195_in_1, msg_to_bit_it_4_vnu_195_in_2, msg_to_bit_it_4_vnu_196_in_0, msg_to_bit_it_4_vnu_196_in_1, msg_to_bit_it_4_vnu_196_in_2, msg_to_bit_it_4_vnu_197_in_0, msg_to_bit_it_4_vnu_197_in_1, msg_to_bit_it_4_vnu_197_in_2, msg_to_bit_it_5_vnu_0_in_0, msg_to_bit_it_5_vnu_0_in_1, msg_to_bit_it_5_vnu_0_in_2, msg_to_bit_it_5_vnu_1_in_0, msg_to_bit_it_5_vnu_1_in_1, msg_to_bit_it_5_vnu_1_in_2, msg_to_bit_it_5_vnu_2_in_0, msg_to_bit_it_5_vnu_2_in_1, msg_to_bit_it_5_vnu_2_in_2, msg_to_bit_it_5_vnu_3_in_0, msg_to_bit_it_5_vnu_3_in_1, msg_to_bit_it_5_vnu_3_in_2, msg_to_bit_it_5_vnu_4_in_0, msg_to_bit_it_5_vnu_4_in_1, msg_to_bit_it_5_vnu_4_in_2, msg_to_bit_it_5_vnu_5_in_0, msg_to_bit_it_5_vnu_5_in_1, msg_to_bit_it_5_vnu_5_in_2, msg_to_bit_it_5_vnu_6_in_0, msg_to_bit_it_5_vnu_6_in_1, msg_to_bit_it_5_vnu_6_in_2, msg_to_bit_it_5_vnu_7_in_0, msg_to_bit_it_5_vnu_7_in_1, msg_to_bit_it_5_vnu_7_in_2, msg_to_bit_it_5_vnu_8_in_0, msg_to_bit_it_5_vnu_8_in_1, msg_to_bit_it_5_vnu_8_in_2, msg_to_bit_it_5_vnu_9_in_0, msg_to_bit_it_5_vnu_9_in_1, msg_to_bit_it_5_vnu_9_in_2, msg_to_bit_it_5_vnu_10_in_0, msg_to_bit_it_5_vnu_10_in_1, msg_to_bit_it_5_vnu_10_in_2, msg_to_bit_it_5_vnu_11_in_0, msg_to_bit_it_5_vnu_11_in_1, msg_to_bit_it_5_vnu_11_in_2, msg_to_bit_it_5_vnu_12_in_0, msg_to_bit_it_5_vnu_12_in_1, msg_to_bit_it_5_vnu_12_in_2, msg_to_bit_it_5_vnu_13_in_0, msg_to_bit_it_5_vnu_13_in_1, msg_to_bit_it_5_vnu_13_in_2, msg_to_bit_it_5_vnu_14_in_0, msg_to_bit_it_5_vnu_14_in_1, msg_to_bit_it_5_vnu_14_in_2, msg_to_bit_it_5_vnu_15_in_0, msg_to_bit_it_5_vnu_15_in_1, msg_to_bit_it_5_vnu_15_in_2, msg_to_bit_it_5_vnu_16_in_0, msg_to_bit_it_5_vnu_16_in_1, msg_to_bit_it_5_vnu_16_in_2, msg_to_bit_it_5_vnu_17_in_0, msg_to_bit_it_5_vnu_17_in_1, msg_to_bit_it_5_vnu_17_in_2, msg_to_bit_it_5_vnu_18_in_0, msg_to_bit_it_5_vnu_18_in_1, msg_to_bit_it_5_vnu_18_in_2, msg_to_bit_it_5_vnu_19_in_0, msg_to_bit_it_5_vnu_19_in_1, msg_to_bit_it_5_vnu_19_in_2, msg_to_bit_it_5_vnu_20_in_0, msg_to_bit_it_5_vnu_20_in_1, msg_to_bit_it_5_vnu_20_in_2, msg_to_bit_it_5_vnu_21_in_0, msg_to_bit_it_5_vnu_21_in_1, msg_to_bit_it_5_vnu_21_in_2, msg_to_bit_it_5_vnu_22_in_0, msg_to_bit_it_5_vnu_22_in_1, msg_to_bit_it_5_vnu_22_in_2, msg_to_bit_it_5_vnu_23_in_0, msg_to_bit_it_5_vnu_23_in_1, msg_to_bit_it_5_vnu_23_in_2, msg_to_bit_it_5_vnu_24_in_0, msg_to_bit_it_5_vnu_24_in_1, msg_to_bit_it_5_vnu_24_in_2, msg_to_bit_it_5_vnu_25_in_0, msg_to_bit_it_5_vnu_25_in_1, msg_to_bit_it_5_vnu_25_in_2, msg_to_bit_it_5_vnu_26_in_0, msg_to_bit_it_5_vnu_26_in_1, msg_to_bit_it_5_vnu_26_in_2, msg_to_bit_it_5_vnu_27_in_0, msg_to_bit_it_5_vnu_27_in_1, msg_to_bit_it_5_vnu_27_in_2, msg_to_bit_it_5_vnu_28_in_0, msg_to_bit_it_5_vnu_28_in_1, msg_to_bit_it_5_vnu_28_in_2, msg_to_bit_it_5_vnu_29_in_0, msg_to_bit_it_5_vnu_29_in_1, msg_to_bit_it_5_vnu_29_in_2, msg_to_bit_it_5_vnu_30_in_0, msg_to_bit_it_5_vnu_30_in_1, msg_to_bit_it_5_vnu_30_in_2, msg_to_bit_it_5_vnu_31_in_0, msg_to_bit_it_5_vnu_31_in_1, msg_to_bit_it_5_vnu_31_in_2, msg_to_bit_it_5_vnu_32_in_0, msg_to_bit_it_5_vnu_32_in_1, msg_to_bit_it_5_vnu_32_in_2, msg_to_bit_it_5_vnu_33_in_0, msg_to_bit_it_5_vnu_33_in_1, msg_to_bit_it_5_vnu_33_in_2, msg_to_bit_it_5_vnu_34_in_0, msg_to_bit_it_5_vnu_34_in_1, msg_to_bit_it_5_vnu_34_in_2, msg_to_bit_it_5_vnu_35_in_0, msg_to_bit_it_5_vnu_35_in_1, msg_to_bit_it_5_vnu_35_in_2, msg_to_bit_it_5_vnu_36_in_0, msg_to_bit_it_5_vnu_36_in_1, msg_to_bit_it_5_vnu_36_in_2, msg_to_bit_it_5_vnu_37_in_0, msg_to_bit_it_5_vnu_37_in_1, msg_to_bit_it_5_vnu_37_in_2, msg_to_bit_it_5_vnu_38_in_0, msg_to_bit_it_5_vnu_38_in_1, msg_to_bit_it_5_vnu_38_in_2, msg_to_bit_it_5_vnu_39_in_0, msg_to_bit_it_5_vnu_39_in_1, msg_to_bit_it_5_vnu_39_in_2, msg_to_bit_it_5_vnu_40_in_0, msg_to_bit_it_5_vnu_40_in_1, msg_to_bit_it_5_vnu_40_in_2, msg_to_bit_it_5_vnu_41_in_0, msg_to_bit_it_5_vnu_41_in_1, msg_to_bit_it_5_vnu_41_in_2, msg_to_bit_it_5_vnu_42_in_0, msg_to_bit_it_5_vnu_42_in_1, msg_to_bit_it_5_vnu_42_in_2, msg_to_bit_it_5_vnu_43_in_0, msg_to_bit_it_5_vnu_43_in_1, msg_to_bit_it_5_vnu_43_in_2, msg_to_bit_it_5_vnu_44_in_0, msg_to_bit_it_5_vnu_44_in_1, msg_to_bit_it_5_vnu_44_in_2, msg_to_bit_it_5_vnu_45_in_0, msg_to_bit_it_5_vnu_45_in_1, msg_to_bit_it_5_vnu_45_in_2, msg_to_bit_it_5_vnu_46_in_0, msg_to_bit_it_5_vnu_46_in_1, msg_to_bit_it_5_vnu_46_in_2, msg_to_bit_it_5_vnu_47_in_0, msg_to_bit_it_5_vnu_47_in_1, msg_to_bit_it_5_vnu_47_in_2, msg_to_bit_it_5_vnu_48_in_0, msg_to_bit_it_5_vnu_48_in_1, msg_to_bit_it_5_vnu_48_in_2, msg_to_bit_it_5_vnu_49_in_0, msg_to_bit_it_5_vnu_49_in_1, msg_to_bit_it_5_vnu_49_in_2, msg_to_bit_it_5_vnu_50_in_0, msg_to_bit_it_5_vnu_50_in_1, msg_to_bit_it_5_vnu_50_in_2, msg_to_bit_it_5_vnu_51_in_0, msg_to_bit_it_5_vnu_51_in_1, msg_to_bit_it_5_vnu_51_in_2, msg_to_bit_it_5_vnu_52_in_0, msg_to_bit_it_5_vnu_52_in_1, msg_to_bit_it_5_vnu_52_in_2, msg_to_bit_it_5_vnu_53_in_0, msg_to_bit_it_5_vnu_53_in_1, msg_to_bit_it_5_vnu_53_in_2, msg_to_bit_it_5_vnu_54_in_0, msg_to_bit_it_5_vnu_54_in_1, msg_to_bit_it_5_vnu_54_in_2, msg_to_bit_it_5_vnu_55_in_0, msg_to_bit_it_5_vnu_55_in_1, msg_to_bit_it_5_vnu_55_in_2, msg_to_bit_it_5_vnu_56_in_0, msg_to_bit_it_5_vnu_56_in_1, msg_to_bit_it_5_vnu_56_in_2, msg_to_bit_it_5_vnu_57_in_0, msg_to_bit_it_5_vnu_57_in_1, msg_to_bit_it_5_vnu_57_in_2, msg_to_bit_it_5_vnu_58_in_0, msg_to_bit_it_5_vnu_58_in_1, msg_to_bit_it_5_vnu_58_in_2, msg_to_bit_it_5_vnu_59_in_0, msg_to_bit_it_5_vnu_59_in_1, msg_to_bit_it_5_vnu_59_in_2, msg_to_bit_it_5_vnu_60_in_0, msg_to_bit_it_5_vnu_60_in_1, msg_to_bit_it_5_vnu_60_in_2, msg_to_bit_it_5_vnu_61_in_0, msg_to_bit_it_5_vnu_61_in_1, msg_to_bit_it_5_vnu_61_in_2, msg_to_bit_it_5_vnu_62_in_0, msg_to_bit_it_5_vnu_62_in_1, msg_to_bit_it_5_vnu_62_in_2, msg_to_bit_it_5_vnu_63_in_0, msg_to_bit_it_5_vnu_63_in_1, msg_to_bit_it_5_vnu_63_in_2, msg_to_bit_it_5_vnu_64_in_0, msg_to_bit_it_5_vnu_64_in_1, msg_to_bit_it_5_vnu_64_in_2, msg_to_bit_it_5_vnu_65_in_0, msg_to_bit_it_5_vnu_65_in_1, msg_to_bit_it_5_vnu_65_in_2, msg_to_bit_it_5_vnu_66_in_0, msg_to_bit_it_5_vnu_66_in_1, msg_to_bit_it_5_vnu_66_in_2, msg_to_bit_it_5_vnu_67_in_0, msg_to_bit_it_5_vnu_67_in_1, msg_to_bit_it_5_vnu_67_in_2, msg_to_bit_it_5_vnu_68_in_0, msg_to_bit_it_5_vnu_68_in_1, msg_to_bit_it_5_vnu_68_in_2, msg_to_bit_it_5_vnu_69_in_0, msg_to_bit_it_5_vnu_69_in_1, msg_to_bit_it_5_vnu_69_in_2, msg_to_bit_it_5_vnu_70_in_0, msg_to_bit_it_5_vnu_70_in_1, msg_to_bit_it_5_vnu_70_in_2, msg_to_bit_it_5_vnu_71_in_0, msg_to_bit_it_5_vnu_71_in_1, msg_to_bit_it_5_vnu_71_in_2, msg_to_bit_it_5_vnu_72_in_0, msg_to_bit_it_5_vnu_72_in_1, msg_to_bit_it_5_vnu_72_in_2, msg_to_bit_it_5_vnu_73_in_0, msg_to_bit_it_5_vnu_73_in_1, msg_to_bit_it_5_vnu_73_in_2, msg_to_bit_it_5_vnu_74_in_0, msg_to_bit_it_5_vnu_74_in_1, msg_to_bit_it_5_vnu_74_in_2, msg_to_bit_it_5_vnu_75_in_0, msg_to_bit_it_5_vnu_75_in_1, msg_to_bit_it_5_vnu_75_in_2, msg_to_bit_it_5_vnu_76_in_0, msg_to_bit_it_5_vnu_76_in_1, msg_to_bit_it_5_vnu_76_in_2, msg_to_bit_it_5_vnu_77_in_0, msg_to_bit_it_5_vnu_77_in_1, msg_to_bit_it_5_vnu_77_in_2, msg_to_bit_it_5_vnu_78_in_0, msg_to_bit_it_5_vnu_78_in_1, msg_to_bit_it_5_vnu_78_in_2, msg_to_bit_it_5_vnu_79_in_0, msg_to_bit_it_5_vnu_79_in_1, msg_to_bit_it_5_vnu_79_in_2, msg_to_bit_it_5_vnu_80_in_0, msg_to_bit_it_5_vnu_80_in_1, msg_to_bit_it_5_vnu_80_in_2, msg_to_bit_it_5_vnu_81_in_0, msg_to_bit_it_5_vnu_81_in_1, msg_to_bit_it_5_vnu_81_in_2, msg_to_bit_it_5_vnu_82_in_0, msg_to_bit_it_5_vnu_82_in_1, msg_to_bit_it_5_vnu_82_in_2, msg_to_bit_it_5_vnu_83_in_0, msg_to_bit_it_5_vnu_83_in_1, msg_to_bit_it_5_vnu_83_in_2, msg_to_bit_it_5_vnu_84_in_0, msg_to_bit_it_5_vnu_84_in_1, msg_to_bit_it_5_vnu_84_in_2, msg_to_bit_it_5_vnu_85_in_0, msg_to_bit_it_5_vnu_85_in_1, msg_to_bit_it_5_vnu_85_in_2, msg_to_bit_it_5_vnu_86_in_0, msg_to_bit_it_5_vnu_86_in_1, msg_to_bit_it_5_vnu_86_in_2, msg_to_bit_it_5_vnu_87_in_0, msg_to_bit_it_5_vnu_87_in_1, msg_to_bit_it_5_vnu_87_in_2, msg_to_bit_it_5_vnu_88_in_0, msg_to_bit_it_5_vnu_88_in_1, msg_to_bit_it_5_vnu_88_in_2, msg_to_bit_it_5_vnu_89_in_0, msg_to_bit_it_5_vnu_89_in_1, msg_to_bit_it_5_vnu_89_in_2, msg_to_bit_it_5_vnu_90_in_0, msg_to_bit_it_5_vnu_90_in_1, msg_to_bit_it_5_vnu_90_in_2, msg_to_bit_it_5_vnu_91_in_0, msg_to_bit_it_5_vnu_91_in_1, msg_to_bit_it_5_vnu_91_in_2, msg_to_bit_it_5_vnu_92_in_0, msg_to_bit_it_5_vnu_92_in_1, msg_to_bit_it_5_vnu_92_in_2, msg_to_bit_it_5_vnu_93_in_0, msg_to_bit_it_5_vnu_93_in_1, msg_to_bit_it_5_vnu_93_in_2, msg_to_bit_it_5_vnu_94_in_0, msg_to_bit_it_5_vnu_94_in_1, msg_to_bit_it_5_vnu_94_in_2, msg_to_bit_it_5_vnu_95_in_0, msg_to_bit_it_5_vnu_95_in_1, msg_to_bit_it_5_vnu_95_in_2, msg_to_bit_it_5_vnu_96_in_0, msg_to_bit_it_5_vnu_96_in_1, msg_to_bit_it_5_vnu_96_in_2, msg_to_bit_it_5_vnu_97_in_0, msg_to_bit_it_5_vnu_97_in_1, msg_to_bit_it_5_vnu_97_in_2, msg_to_bit_it_5_vnu_98_in_0, msg_to_bit_it_5_vnu_98_in_1, msg_to_bit_it_5_vnu_98_in_2, msg_to_bit_it_5_vnu_99_in_0, msg_to_bit_it_5_vnu_99_in_1, msg_to_bit_it_5_vnu_99_in_2, msg_to_bit_it_5_vnu_100_in_0, msg_to_bit_it_5_vnu_100_in_1, msg_to_bit_it_5_vnu_100_in_2, msg_to_bit_it_5_vnu_101_in_0, msg_to_bit_it_5_vnu_101_in_1, msg_to_bit_it_5_vnu_101_in_2, msg_to_bit_it_5_vnu_102_in_0, msg_to_bit_it_5_vnu_102_in_1, msg_to_bit_it_5_vnu_102_in_2, msg_to_bit_it_5_vnu_103_in_0, msg_to_bit_it_5_vnu_103_in_1, msg_to_bit_it_5_vnu_103_in_2, msg_to_bit_it_5_vnu_104_in_0, msg_to_bit_it_5_vnu_104_in_1, msg_to_bit_it_5_vnu_104_in_2, msg_to_bit_it_5_vnu_105_in_0, msg_to_bit_it_5_vnu_105_in_1, msg_to_bit_it_5_vnu_105_in_2, msg_to_bit_it_5_vnu_106_in_0, msg_to_bit_it_5_vnu_106_in_1, msg_to_bit_it_5_vnu_106_in_2, msg_to_bit_it_5_vnu_107_in_0, msg_to_bit_it_5_vnu_107_in_1, msg_to_bit_it_5_vnu_107_in_2, msg_to_bit_it_5_vnu_108_in_0, msg_to_bit_it_5_vnu_108_in_1, msg_to_bit_it_5_vnu_108_in_2, msg_to_bit_it_5_vnu_109_in_0, msg_to_bit_it_5_vnu_109_in_1, msg_to_bit_it_5_vnu_109_in_2, msg_to_bit_it_5_vnu_110_in_0, msg_to_bit_it_5_vnu_110_in_1, msg_to_bit_it_5_vnu_110_in_2, msg_to_bit_it_5_vnu_111_in_0, msg_to_bit_it_5_vnu_111_in_1, msg_to_bit_it_5_vnu_111_in_2, msg_to_bit_it_5_vnu_112_in_0, msg_to_bit_it_5_vnu_112_in_1, msg_to_bit_it_5_vnu_112_in_2, msg_to_bit_it_5_vnu_113_in_0, msg_to_bit_it_5_vnu_113_in_1, msg_to_bit_it_5_vnu_113_in_2, msg_to_bit_it_5_vnu_114_in_0, msg_to_bit_it_5_vnu_114_in_1, msg_to_bit_it_5_vnu_114_in_2, msg_to_bit_it_5_vnu_115_in_0, msg_to_bit_it_5_vnu_115_in_1, msg_to_bit_it_5_vnu_115_in_2, msg_to_bit_it_5_vnu_116_in_0, msg_to_bit_it_5_vnu_116_in_1, msg_to_bit_it_5_vnu_116_in_2, msg_to_bit_it_5_vnu_117_in_0, msg_to_bit_it_5_vnu_117_in_1, msg_to_bit_it_5_vnu_117_in_2, msg_to_bit_it_5_vnu_118_in_0, msg_to_bit_it_5_vnu_118_in_1, msg_to_bit_it_5_vnu_118_in_2, msg_to_bit_it_5_vnu_119_in_0, msg_to_bit_it_5_vnu_119_in_1, msg_to_bit_it_5_vnu_119_in_2, msg_to_bit_it_5_vnu_120_in_0, msg_to_bit_it_5_vnu_120_in_1, msg_to_bit_it_5_vnu_120_in_2, msg_to_bit_it_5_vnu_121_in_0, msg_to_bit_it_5_vnu_121_in_1, msg_to_bit_it_5_vnu_121_in_2, msg_to_bit_it_5_vnu_122_in_0, msg_to_bit_it_5_vnu_122_in_1, msg_to_bit_it_5_vnu_122_in_2, msg_to_bit_it_5_vnu_123_in_0, msg_to_bit_it_5_vnu_123_in_1, msg_to_bit_it_5_vnu_123_in_2, msg_to_bit_it_5_vnu_124_in_0, msg_to_bit_it_5_vnu_124_in_1, msg_to_bit_it_5_vnu_124_in_2, msg_to_bit_it_5_vnu_125_in_0, msg_to_bit_it_5_vnu_125_in_1, msg_to_bit_it_5_vnu_125_in_2, msg_to_bit_it_5_vnu_126_in_0, msg_to_bit_it_5_vnu_126_in_1, msg_to_bit_it_5_vnu_126_in_2, msg_to_bit_it_5_vnu_127_in_0, msg_to_bit_it_5_vnu_127_in_1, msg_to_bit_it_5_vnu_127_in_2, msg_to_bit_it_5_vnu_128_in_0, msg_to_bit_it_5_vnu_128_in_1, msg_to_bit_it_5_vnu_128_in_2, msg_to_bit_it_5_vnu_129_in_0, msg_to_bit_it_5_vnu_129_in_1, msg_to_bit_it_5_vnu_129_in_2, msg_to_bit_it_5_vnu_130_in_0, msg_to_bit_it_5_vnu_130_in_1, msg_to_bit_it_5_vnu_130_in_2, msg_to_bit_it_5_vnu_131_in_0, msg_to_bit_it_5_vnu_131_in_1, msg_to_bit_it_5_vnu_131_in_2, msg_to_bit_it_5_vnu_132_in_0, msg_to_bit_it_5_vnu_132_in_1, msg_to_bit_it_5_vnu_132_in_2, msg_to_bit_it_5_vnu_133_in_0, msg_to_bit_it_5_vnu_133_in_1, msg_to_bit_it_5_vnu_133_in_2, msg_to_bit_it_5_vnu_134_in_0, msg_to_bit_it_5_vnu_134_in_1, msg_to_bit_it_5_vnu_134_in_2, msg_to_bit_it_5_vnu_135_in_0, msg_to_bit_it_5_vnu_135_in_1, msg_to_bit_it_5_vnu_135_in_2, msg_to_bit_it_5_vnu_136_in_0, msg_to_bit_it_5_vnu_136_in_1, msg_to_bit_it_5_vnu_136_in_2, msg_to_bit_it_5_vnu_137_in_0, msg_to_bit_it_5_vnu_137_in_1, msg_to_bit_it_5_vnu_137_in_2, msg_to_bit_it_5_vnu_138_in_0, msg_to_bit_it_5_vnu_138_in_1, msg_to_bit_it_5_vnu_138_in_2, msg_to_bit_it_5_vnu_139_in_0, msg_to_bit_it_5_vnu_139_in_1, msg_to_bit_it_5_vnu_139_in_2, msg_to_bit_it_5_vnu_140_in_0, msg_to_bit_it_5_vnu_140_in_1, msg_to_bit_it_5_vnu_140_in_2, msg_to_bit_it_5_vnu_141_in_0, msg_to_bit_it_5_vnu_141_in_1, msg_to_bit_it_5_vnu_141_in_2, msg_to_bit_it_5_vnu_142_in_0, msg_to_bit_it_5_vnu_142_in_1, msg_to_bit_it_5_vnu_142_in_2, msg_to_bit_it_5_vnu_143_in_0, msg_to_bit_it_5_vnu_143_in_1, msg_to_bit_it_5_vnu_143_in_2, msg_to_bit_it_5_vnu_144_in_0, msg_to_bit_it_5_vnu_144_in_1, msg_to_bit_it_5_vnu_144_in_2, msg_to_bit_it_5_vnu_145_in_0, msg_to_bit_it_5_vnu_145_in_1, msg_to_bit_it_5_vnu_145_in_2, msg_to_bit_it_5_vnu_146_in_0, msg_to_bit_it_5_vnu_146_in_1, msg_to_bit_it_5_vnu_146_in_2, msg_to_bit_it_5_vnu_147_in_0, msg_to_bit_it_5_vnu_147_in_1, msg_to_bit_it_5_vnu_147_in_2, msg_to_bit_it_5_vnu_148_in_0, msg_to_bit_it_5_vnu_148_in_1, msg_to_bit_it_5_vnu_148_in_2, msg_to_bit_it_5_vnu_149_in_0, msg_to_bit_it_5_vnu_149_in_1, msg_to_bit_it_5_vnu_149_in_2, msg_to_bit_it_5_vnu_150_in_0, msg_to_bit_it_5_vnu_150_in_1, msg_to_bit_it_5_vnu_150_in_2, msg_to_bit_it_5_vnu_151_in_0, msg_to_bit_it_5_vnu_151_in_1, msg_to_bit_it_5_vnu_151_in_2, msg_to_bit_it_5_vnu_152_in_0, msg_to_bit_it_5_vnu_152_in_1, msg_to_bit_it_5_vnu_152_in_2, msg_to_bit_it_5_vnu_153_in_0, msg_to_bit_it_5_vnu_153_in_1, msg_to_bit_it_5_vnu_153_in_2, msg_to_bit_it_5_vnu_154_in_0, msg_to_bit_it_5_vnu_154_in_1, msg_to_bit_it_5_vnu_154_in_2, msg_to_bit_it_5_vnu_155_in_0, msg_to_bit_it_5_vnu_155_in_1, msg_to_bit_it_5_vnu_155_in_2, msg_to_bit_it_5_vnu_156_in_0, msg_to_bit_it_5_vnu_156_in_1, msg_to_bit_it_5_vnu_156_in_2, msg_to_bit_it_5_vnu_157_in_0, msg_to_bit_it_5_vnu_157_in_1, msg_to_bit_it_5_vnu_157_in_2, msg_to_bit_it_5_vnu_158_in_0, msg_to_bit_it_5_vnu_158_in_1, msg_to_bit_it_5_vnu_158_in_2, msg_to_bit_it_5_vnu_159_in_0, msg_to_bit_it_5_vnu_159_in_1, msg_to_bit_it_5_vnu_159_in_2, msg_to_bit_it_5_vnu_160_in_0, msg_to_bit_it_5_vnu_160_in_1, msg_to_bit_it_5_vnu_160_in_2, msg_to_bit_it_5_vnu_161_in_0, msg_to_bit_it_5_vnu_161_in_1, msg_to_bit_it_5_vnu_161_in_2, msg_to_bit_it_5_vnu_162_in_0, msg_to_bit_it_5_vnu_162_in_1, msg_to_bit_it_5_vnu_162_in_2, msg_to_bit_it_5_vnu_163_in_0, msg_to_bit_it_5_vnu_163_in_1, msg_to_bit_it_5_vnu_163_in_2, msg_to_bit_it_5_vnu_164_in_0, msg_to_bit_it_5_vnu_164_in_1, msg_to_bit_it_5_vnu_164_in_2, msg_to_bit_it_5_vnu_165_in_0, msg_to_bit_it_5_vnu_165_in_1, msg_to_bit_it_5_vnu_165_in_2, msg_to_bit_it_5_vnu_166_in_0, msg_to_bit_it_5_vnu_166_in_1, msg_to_bit_it_5_vnu_166_in_2, msg_to_bit_it_5_vnu_167_in_0, msg_to_bit_it_5_vnu_167_in_1, msg_to_bit_it_5_vnu_167_in_2, msg_to_bit_it_5_vnu_168_in_0, msg_to_bit_it_5_vnu_168_in_1, msg_to_bit_it_5_vnu_168_in_2, msg_to_bit_it_5_vnu_169_in_0, msg_to_bit_it_5_vnu_169_in_1, msg_to_bit_it_5_vnu_169_in_2, msg_to_bit_it_5_vnu_170_in_0, msg_to_bit_it_5_vnu_170_in_1, msg_to_bit_it_5_vnu_170_in_2, msg_to_bit_it_5_vnu_171_in_0, msg_to_bit_it_5_vnu_171_in_1, msg_to_bit_it_5_vnu_171_in_2, msg_to_bit_it_5_vnu_172_in_0, msg_to_bit_it_5_vnu_172_in_1, msg_to_bit_it_5_vnu_172_in_2, msg_to_bit_it_5_vnu_173_in_0, msg_to_bit_it_5_vnu_173_in_1, msg_to_bit_it_5_vnu_173_in_2, msg_to_bit_it_5_vnu_174_in_0, msg_to_bit_it_5_vnu_174_in_1, msg_to_bit_it_5_vnu_174_in_2, msg_to_bit_it_5_vnu_175_in_0, msg_to_bit_it_5_vnu_175_in_1, msg_to_bit_it_5_vnu_175_in_2, msg_to_bit_it_5_vnu_176_in_0, msg_to_bit_it_5_vnu_176_in_1, msg_to_bit_it_5_vnu_176_in_2, msg_to_bit_it_5_vnu_177_in_0, msg_to_bit_it_5_vnu_177_in_1, msg_to_bit_it_5_vnu_177_in_2, msg_to_bit_it_5_vnu_178_in_0, msg_to_bit_it_5_vnu_178_in_1, msg_to_bit_it_5_vnu_178_in_2, msg_to_bit_it_5_vnu_179_in_0, msg_to_bit_it_5_vnu_179_in_1, msg_to_bit_it_5_vnu_179_in_2, msg_to_bit_it_5_vnu_180_in_0, msg_to_bit_it_5_vnu_180_in_1, msg_to_bit_it_5_vnu_180_in_2, msg_to_bit_it_5_vnu_181_in_0, msg_to_bit_it_5_vnu_181_in_1, msg_to_bit_it_5_vnu_181_in_2, msg_to_bit_it_5_vnu_182_in_0, msg_to_bit_it_5_vnu_182_in_1, msg_to_bit_it_5_vnu_182_in_2, msg_to_bit_it_5_vnu_183_in_0, msg_to_bit_it_5_vnu_183_in_1, msg_to_bit_it_5_vnu_183_in_2, msg_to_bit_it_5_vnu_184_in_0, msg_to_bit_it_5_vnu_184_in_1, msg_to_bit_it_5_vnu_184_in_2, msg_to_bit_it_5_vnu_185_in_0, msg_to_bit_it_5_vnu_185_in_1, msg_to_bit_it_5_vnu_185_in_2, msg_to_bit_it_5_vnu_186_in_0, msg_to_bit_it_5_vnu_186_in_1, msg_to_bit_it_5_vnu_186_in_2, msg_to_bit_it_5_vnu_187_in_0, msg_to_bit_it_5_vnu_187_in_1, msg_to_bit_it_5_vnu_187_in_2, msg_to_bit_it_5_vnu_188_in_0, msg_to_bit_it_5_vnu_188_in_1, msg_to_bit_it_5_vnu_188_in_2, msg_to_bit_it_5_vnu_189_in_0, msg_to_bit_it_5_vnu_189_in_1, msg_to_bit_it_5_vnu_189_in_2, msg_to_bit_it_5_vnu_190_in_0, msg_to_bit_it_5_vnu_190_in_1, msg_to_bit_it_5_vnu_190_in_2, msg_to_bit_it_5_vnu_191_in_0, msg_to_bit_it_5_vnu_191_in_1, msg_to_bit_it_5_vnu_191_in_2, msg_to_bit_it_5_vnu_192_in_0, msg_to_bit_it_5_vnu_192_in_1, msg_to_bit_it_5_vnu_192_in_2, msg_to_bit_it_5_vnu_193_in_0, msg_to_bit_it_5_vnu_193_in_1, msg_to_bit_it_5_vnu_193_in_2, msg_to_bit_it_5_vnu_194_in_0, msg_to_bit_it_5_vnu_194_in_1, msg_to_bit_it_5_vnu_194_in_2, msg_to_bit_it_5_vnu_195_in_0, msg_to_bit_it_5_vnu_195_in_1, msg_to_bit_it_5_vnu_195_in_2, msg_to_bit_it_5_vnu_196_in_0, msg_to_bit_it_5_vnu_196_in_1, msg_to_bit_it_5_vnu_196_in_2, msg_to_bit_it_5_vnu_197_in_0, msg_to_bit_it_5_vnu_197_in_1, msg_to_bit_it_5_vnu_197_in_2, msg_to_bit_it_6_vnu_0_in_0, msg_to_bit_it_6_vnu_0_in_1, msg_to_bit_it_6_vnu_0_in_2, msg_to_bit_it_6_vnu_1_in_0, msg_to_bit_it_6_vnu_1_in_1, msg_to_bit_it_6_vnu_1_in_2, msg_to_bit_it_6_vnu_2_in_0, msg_to_bit_it_6_vnu_2_in_1, msg_to_bit_it_6_vnu_2_in_2, msg_to_bit_it_6_vnu_3_in_0, msg_to_bit_it_6_vnu_3_in_1, msg_to_bit_it_6_vnu_3_in_2, msg_to_bit_it_6_vnu_4_in_0, msg_to_bit_it_6_vnu_4_in_1, msg_to_bit_it_6_vnu_4_in_2, msg_to_bit_it_6_vnu_5_in_0, msg_to_bit_it_6_vnu_5_in_1, msg_to_bit_it_6_vnu_5_in_2, msg_to_bit_it_6_vnu_6_in_0, msg_to_bit_it_6_vnu_6_in_1, msg_to_bit_it_6_vnu_6_in_2, msg_to_bit_it_6_vnu_7_in_0, msg_to_bit_it_6_vnu_7_in_1, msg_to_bit_it_6_vnu_7_in_2, msg_to_bit_it_6_vnu_8_in_0, msg_to_bit_it_6_vnu_8_in_1, msg_to_bit_it_6_vnu_8_in_2, msg_to_bit_it_6_vnu_9_in_0, msg_to_bit_it_6_vnu_9_in_1, msg_to_bit_it_6_vnu_9_in_2, msg_to_bit_it_6_vnu_10_in_0, msg_to_bit_it_6_vnu_10_in_1, msg_to_bit_it_6_vnu_10_in_2, msg_to_bit_it_6_vnu_11_in_0, msg_to_bit_it_6_vnu_11_in_1, msg_to_bit_it_6_vnu_11_in_2, msg_to_bit_it_6_vnu_12_in_0, msg_to_bit_it_6_vnu_12_in_1, msg_to_bit_it_6_vnu_12_in_2, msg_to_bit_it_6_vnu_13_in_0, msg_to_bit_it_6_vnu_13_in_1, msg_to_bit_it_6_vnu_13_in_2, msg_to_bit_it_6_vnu_14_in_0, msg_to_bit_it_6_vnu_14_in_1, msg_to_bit_it_6_vnu_14_in_2, msg_to_bit_it_6_vnu_15_in_0, msg_to_bit_it_6_vnu_15_in_1, msg_to_bit_it_6_vnu_15_in_2, msg_to_bit_it_6_vnu_16_in_0, msg_to_bit_it_6_vnu_16_in_1, msg_to_bit_it_6_vnu_16_in_2, msg_to_bit_it_6_vnu_17_in_0, msg_to_bit_it_6_vnu_17_in_1, msg_to_bit_it_6_vnu_17_in_2, msg_to_bit_it_6_vnu_18_in_0, msg_to_bit_it_6_vnu_18_in_1, msg_to_bit_it_6_vnu_18_in_2, msg_to_bit_it_6_vnu_19_in_0, msg_to_bit_it_6_vnu_19_in_1, msg_to_bit_it_6_vnu_19_in_2, msg_to_bit_it_6_vnu_20_in_0, msg_to_bit_it_6_vnu_20_in_1, msg_to_bit_it_6_vnu_20_in_2, msg_to_bit_it_6_vnu_21_in_0, msg_to_bit_it_6_vnu_21_in_1, msg_to_bit_it_6_vnu_21_in_2, msg_to_bit_it_6_vnu_22_in_0, msg_to_bit_it_6_vnu_22_in_1, msg_to_bit_it_6_vnu_22_in_2, msg_to_bit_it_6_vnu_23_in_0, msg_to_bit_it_6_vnu_23_in_1, msg_to_bit_it_6_vnu_23_in_2, msg_to_bit_it_6_vnu_24_in_0, msg_to_bit_it_6_vnu_24_in_1, msg_to_bit_it_6_vnu_24_in_2, msg_to_bit_it_6_vnu_25_in_0, msg_to_bit_it_6_vnu_25_in_1, msg_to_bit_it_6_vnu_25_in_2, msg_to_bit_it_6_vnu_26_in_0, msg_to_bit_it_6_vnu_26_in_1, msg_to_bit_it_6_vnu_26_in_2, msg_to_bit_it_6_vnu_27_in_0, msg_to_bit_it_6_vnu_27_in_1, msg_to_bit_it_6_vnu_27_in_2, msg_to_bit_it_6_vnu_28_in_0, msg_to_bit_it_6_vnu_28_in_1, msg_to_bit_it_6_vnu_28_in_2, msg_to_bit_it_6_vnu_29_in_0, msg_to_bit_it_6_vnu_29_in_1, msg_to_bit_it_6_vnu_29_in_2, msg_to_bit_it_6_vnu_30_in_0, msg_to_bit_it_6_vnu_30_in_1, msg_to_bit_it_6_vnu_30_in_2, msg_to_bit_it_6_vnu_31_in_0, msg_to_bit_it_6_vnu_31_in_1, msg_to_bit_it_6_vnu_31_in_2, msg_to_bit_it_6_vnu_32_in_0, msg_to_bit_it_6_vnu_32_in_1, msg_to_bit_it_6_vnu_32_in_2, msg_to_bit_it_6_vnu_33_in_0, msg_to_bit_it_6_vnu_33_in_1, msg_to_bit_it_6_vnu_33_in_2, msg_to_bit_it_6_vnu_34_in_0, msg_to_bit_it_6_vnu_34_in_1, msg_to_bit_it_6_vnu_34_in_2, msg_to_bit_it_6_vnu_35_in_0, msg_to_bit_it_6_vnu_35_in_1, msg_to_bit_it_6_vnu_35_in_2, msg_to_bit_it_6_vnu_36_in_0, msg_to_bit_it_6_vnu_36_in_1, msg_to_bit_it_6_vnu_36_in_2, msg_to_bit_it_6_vnu_37_in_0, msg_to_bit_it_6_vnu_37_in_1, msg_to_bit_it_6_vnu_37_in_2, msg_to_bit_it_6_vnu_38_in_0, msg_to_bit_it_6_vnu_38_in_1, msg_to_bit_it_6_vnu_38_in_2, msg_to_bit_it_6_vnu_39_in_0, msg_to_bit_it_6_vnu_39_in_1, msg_to_bit_it_6_vnu_39_in_2, msg_to_bit_it_6_vnu_40_in_0, msg_to_bit_it_6_vnu_40_in_1, msg_to_bit_it_6_vnu_40_in_2, msg_to_bit_it_6_vnu_41_in_0, msg_to_bit_it_6_vnu_41_in_1, msg_to_bit_it_6_vnu_41_in_2, msg_to_bit_it_6_vnu_42_in_0, msg_to_bit_it_6_vnu_42_in_1, msg_to_bit_it_6_vnu_42_in_2, msg_to_bit_it_6_vnu_43_in_0, msg_to_bit_it_6_vnu_43_in_1, msg_to_bit_it_6_vnu_43_in_2, msg_to_bit_it_6_vnu_44_in_0, msg_to_bit_it_6_vnu_44_in_1, msg_to_bit_it_6_vnu_44_in_2, msg_to_bit_it_6_vnu_45_in_0, msg_to_bit_it_6_vnu_45_in_1, msg_to_bit_it_6_vnu_45_in_2, msg_to_bit_it_6_vnu_46_in_0, msg_to_bit_it_6_vnu_46_in_1, msg_to_bit_it_6_vnu_46_in_2, msg_to_bit_it_6_vnu_47_in_0, msg_to_bit_it_6_vnu_47_in_1, msg_to_bit_it_6_vnu_47_in_2, msg_to_bit_it_6_vnu_48_in_0, msg_to_bit_it_6_vnu_48_in_1, msg_to_bit_it_6_vnu_48_in_2, msg_to_bit_it_6_vnu_49_in_0, msg_to_bit_it_6_vnu_49_in_1, msg_to_bit_it_6_vnu_49_in_2, msg_to_bit_it_6_vnu_50_in_0, msg_to_bit_it_6_vnu_50_in_1, msg_to_bit_it_6_vnu_50_in_2, msg_to_bit_it_6_vnu_51_in_0, msg_to_bit_it_6_vnu_51_in_1, msg_to_bit_it_6_vnu_51_in_2, msg_to_bit_it_6_vnu_52_in_0, msg_to_bit_it_6_vnu_52_in_1, msg_to_bit_it_6_vnu_52_in_2, msg_to_bit_it_6_vnu_53_in_0, msg_to_bit_it_6_vnu_53_in_1, msg_to_bit_it_6_vnu_53_in_2, msg_to_bit_it_6_vnu_54_in_0, msg_to_bit_it_6_vnu_54_in_1, msg_to_bit_it_6_vnu_54_in_2, msg_to_bit_it_6_vnu_55_in_0, msg_to_bit_it_6_vnu_55_in_1, msg_to_bit_it_6_vnu_55_in_2, msg_to_bit_it_6_vnu_56_in_0, msg_to_bit_it_6_vnu_56_in_1, msg_to_bit_it_6_vnu_56_in_2, msg_to_bit_it_6_vnu_57_in_0, msg_to_bit_it_6_vnu_57_in_1, msg_to_bit_it_6_vnu_57_in_2, msg_to_bit_it_6_vnu_58_in_0, msg_to_bit_it_6_vnu_58_in_1, msg_to_bit_it_6_vnu_58_in_2, msg_to_bit_it_6_vnu_59_in_0, msg_to_bit_it_6_vnu_59_in_1, msg_to_bit_it_6_vnu_59_in_2, msg_to_bit_it_6_vnu_60_in_0, msg_to_bit_it_6_vnu_60_in_1, msg_to_bit_it_6_vnu_60_in_2, msg_to_bit_it_6_vnu_61_in_0, msg_to_bit_it_6_vnu_61_in_1, msg_to_bit_it_6_vnu_61_in_2, msg_to_bit_it_6_vnu_62_in_0, msg_to_bit_it_6_vnu_62_in_1, msg_to_bit_it_6_vnu_62_in_2, msg_to_bit_it_6_vnu_63_in_0, msg_to_bit_it_6_vnu_63_in_1, msg_to_bit_it_6_vnu_63_in_2, msg_to_bit_it_6_vnu_64_in_0, msg_to_bit_it_6_vnu_64_in_1, msg_to_bit_it_6_vnu_64_in_2, msg_to_bit_it_6_vnu_65_in_0, msg_to_bit_it_6_vnu_65_in_1, msg_to_bit_it_6_vnu_65_in_2, msg_to_bit_it_6_vnu_66_in_0, msg_to_bit_it_6_vnu_66_in_1, msg_to_bit_it_6_vnu_66_in_2, msg_to_bit_it_6_vnu_67_in_0, msg_to_bit_it_6_vnu_67_in_1, msg_to_bit_it_6_vnu_67_in_2, msg_to_bit_it_6_vnu_68_in_0, msg_to_bit_it_6_vnu_68_in_1, msg_to_bit_it_6_vnu_68_in_2, msg_to_bit_it_6_vnu_69_in_0, msg_to_bit_it_6_vnu_69_in_1, msg_to_bit_it_6_vnu_69_in_2, msg_to_bit_it_6_vnu_70_in_0, msg_to_bit_it_6_vnu_70_in_1, msg_to_bit_it_6_vnu_70_in_2, msg_to_bit_it_6_vnu_71_in_0, msg_to_bit_it_6_vnu_71_in_1, msg_to_bit_it_6_vnu_71_in_2, msg_to_bit_it_6_vnu_72_in_0, msg_to_bit_it_6_vnu_72_in_1, msg_to_bit_it_6_vnu_72_in_2, msg_to_bit_it_6_vnu_73_in_0, msg_to_bit_it_6_vnu_73_in_1, msg_to_bit_it_6_vnu_73_in_2, msg_to_bit_it_6_vnu_74_in_0, msg_to_bit_it_6_vnu_74_in_1, msg_to_bit_it_6_vnu_74_in_2, msg_to_bit_it_6_vnu_75_in_0, msg_to_bit_it_6_vnu_75_in_1, msg_to_bit_it_6_vnu_75_in_2, msg_to_bit_it_6_vnu_76_in_0, msg_to_bit_it_6_vnu_76_in_1, msg_to_bit_it_6_vnu_76_in_2, msg_to_bit_it_6_vnu_77_in_0, msg_to_bit_it_6_vnu_77_in_1, msg_to_bit_it_6_vnu_77_in_2, msg_to_bit_it_6_vnu_78_in_0, msg_to_bit_it_6_vnu_78_in_1, msg_to_bit_it_6_vnu_78_in_2, msg_to_bit_it_6_vnu_79_in_0, msg_to_bit_it_6_vnu_79_in_1, msg_to_bit_it_6_vnu_79_in_2, msg_to_bit_it_6_vnu_80_in_0, msg_to_bit_it_6_vnu_80_in_1, msg_to_bit_it_6_vnu_80_in_2, msg_to_bit_it_6_vnu_81_in_0, msg_to_bit_it_6_vnu_81_in_1, msg_to_bit_it_6_vnu_81_in_2, msg_to_bit_it_6_vnu_82_in_0, msg_to_bit_it_6_vnu_82_in_1, msg_to_bit_it_6_vnu_82_in_2, msg_to_bit_it_6_vnu_83_in_0, msg_to_bit_it_6_vnu_83_in_1, msg_to_bit_it_6_vnu_83_in_2, msg_to_bit_it_6_vnu_84_in_0, msg_to_bit_it_6_vnu_84_in_1, msg_to_bit_it_6_vnu_84_in_2, msg_to_bit_it_6_vnu_85_in_0, msg_to_bit_it_6_vnu_85_in_1, msg_to_bit_it_6_vnu_85_in_2, msg_to_bit_it_6_vnu_86_in_0, msg_to_bit_it_6_vnu_86_in_1, msg_to_bit_it_6_vnu_86_in_2, msg_to_bit_it_6_vnu_87_in_0, msg_to_bit_it_6_vnu_87_in_1, msg_to_bit_it_6_vnu_87_in_2, msg_to_bit_it_6_vnu_88_in_0, msg_to_bit_it_6_vnu_88_in_1, msg_to_bit_it_6_vnu_88_in_2, msg_to_bit_it_6_vnu_89_in_0, msg_to_bit_it_6_vnu_89_in_1, msg_to_bit_it_6_vnu_89_in_2, msg_to_bit_it_6_vnu_90_in_0, msg_to_bit_it_6_vnu_90_in_1, msg_to_bit_it_6_vnu_90_in_2, msg_to_bit_it_6_vnu_91_in_0, msg_to_bit_it_6_vnu_91_in_1, msg_to_bit_it_6_vnu_91_in_2, msg_to_bit_it_6_vnu_92_in_0, msg_to_bit_it_6_vnu_92_in_1, msg_to_bit_it_6_vnu_92_in_2, msg_to_bit_it_6_vnu_93_in_0, msg_to_bit_it_6_vnu_93_in_1, msg_to_bit_it_6_vnu_93_in_2, msg_to_bit_it_6_vnu_94_in_0, msg_to_bit_it_6_vnu_94_in_1, msg_to_bit_it_6_vnu_94_in_2, msg_to_bit_it_6_vnu_95_in_0, msg_to_bit_it_6_vnu_95_in_1, msg_to_bit_it_6_vnu_95_in_2, msg_to_bit_it_6_vnu_96_in_0, msg_to_bit_it_6_vnu_96_in_1, msg_to_bit_it_6_vnu_96_in_2, msg_to_bit_it_6_vnu_97_in_0, msg_to_bit_it_6_vnu_97_in_1, msg_to_bit_it_6_vnu_97_in_2, msg_to_bit_it_6_vnu_98_in_0, msg_to_bit_it_6_vnu_98_in_1, msg_to_bit_it_6_vnu_98_in_2, msg_to_bit_it_6_vnu_99_in_0, msg_to_bit_it_6_vnu_99_in_1, msg_to_bit_it_6_vnu_99_in_2, msg_to_bit_it_6_vnu_100_in_0, msg_to_bit_it_6_vnu_100_in_1, msg_to_bit_it_6_vnu_100_in_2, msg_to_bit_it_6_vnu_101_in_0, msg_to_bit_it_6_vnu_101_in_1, msg_to_bit_it_6_vnu_101_in_2, msg_to_bit_it_6_vnu_102_in_0, msg_to_bit_it_6_vnu_102_in_1, msg_to_bit_it_6_vnu_102_in_2, msg_to_bit_it_6_vnu_103_in_0, msg_to_bit_it_6_vnu_103_in_1, msg_to_bit_it_6_vnu_103_in_2, msg_to_bit_it_6_vnu_104_in_0, msg_to_bit_it_6_vnu_104_in_1, msg_to_bit_it_6_vnu_104_in_2, msg_to_bit_it_6_vnu_105_in_0, msg_to_bit_it_6_vnu_105_in_1, msg_to_bit_it_6_vnu_105_in_2, msg_to_bit_it_6_vnu_106_in_0, msg_to_bit_it_6_vnu_106_in_1, msg_to_bit_it_6_vnu_106_in_2, msg_to_bit_it_6_vnu_107_in_0, msg_to_bit_it_6_vnu_107_in_1, msg_to_bit_it_6_vnu_107_in_2, msg_to_bit_it_6_vnu_108_in_0, msg_to_bit_it_6_vnu_108_in_1, msg_to_bit_it_6_vnu_108_in_2, msg_to_bit_it_6_vnu_109_in_0, msg_to_bit_it_6_vnu_109_in_1, msg_to_bit_it_6_vnu_109_in_2, msg_to_bit_it_6_vnu_110_in_0, msg_to_bit_it_6_vnu_110_in_1, msg_to_bit_it_6_vnu_110_in_2, msg_to_bit_it_6_vnu_111_in_0, msg_to_bit_it_6_vnu_111_in_1, msg_to_bit_it_6_vnu_111_in_2, msg_to_bit_it_6_vnu_112_in_0, msg_to_bit_it_6_vnu_112_in_1, msg_to_bit_it_6_vnu_112_in_2, msg_to_bit_it_6_vnu_113_in_0, msg_to_bit_it_6_vnu_113_in_1, msg_to_bit_it_6_vnu_113_in_2, msg_to_bit_it_6_vnu_114_in_0, msg_to_bit_it_6_vnu_114_in_1, msg_to_bit_it_6_vnu_114_in_2, msg_to_bit_it_6_vnu_115_in_0, msg_to_bit_it_6_vnu_115_in_1, msg_to_bit_it_6_vnu_115_in_2, msg_to_bit_it_6_vnu_116_in_0, msg_to_bit_it_6_vnu_116_in_1, msg_to_bit_it_6_vnu_116_in_2, msg_to_bit_it_6_vnu_117_in_0, msg_to_bit_it_6_vnu_117_in_1, msg_to_bit_it_6_vnu_117_in_2, msg_to_bit_it_6_vnu_118_in_0, msg_to_bit_it_6_vnu_118_in_1, msg_to_bit_it_6_vnu_118_in_2, msg_to_bit_it_6_vnu_119_in_0, msg_to_bit_it_6_vnu_119_in_1, msg_to_bit_it_6_vnu_119_in_2, msg_to_bit_it_6_vnu_120_in_0, msg_to_bit_it_6_vnu_120_in_1, msg_to_bit_it_6_vnu_120_in_2, msg_to_bit_it_6_vnu_121_in_0, msg_to_bit_it_6_vnu_121_in_1, msg_to_bit_it_6_vnu_121_in_2, msg_to_bit_it_6_vnu_122_in_0, msg_to_bit_it_6_vnu_122_in_1, msg_to_bit_it_6_vnu_122_in_2, msg_to_bit_it_6_vnu_123_in_0, msg_to_bit_it_6_vnu_123_in_1, msg_to_bit_it_6_vnu_123_in_2, msg_to_bit_it_6_vnu_124_in_0, msg_to_bit_it_6_vnu_124_in_1, msg_to_bit_it_6_vnu_124_in_2, msg_to_bit_it_6_vnu_125_in_0, msg_to_bit_it_6_vnu_125_in_1, msg_to_bit_it_6_vnu_125_in_2, msg_to_bit_it_6_vnu_126_in_0, msg_to_bit_it_6_vnu_126_in_1, msg_to_bit_it_6_vnu_126_in_2, msg_to_bit_it_6_vnu_127_in_0, msg_to_bit_it_6_vnu_127_in_1, msg_to_bit_it_6_vnu_127_in_2, msg_to_bit_it_6_vnu_128_in_0, msg_to_bit_it_6_vnu_128_in_1, msg_to_bit_it_6_vnu_128_in_2, msg_to_bit_it_6_vnu_129_in_0, msg_to_bit_it_6_vnu_129_in_1, msg_to_bit_it_6_vnu_129_in_2, msg_to_bit_it_6_vnu_130_in_0, msg_to_bit_it_6_vnu_130_in_1, msg_to_bit_it_6_vnu_130_in_2, msg_to_bit_it_6_vnu_131_in_0, msg_to_bit_it_6_vnu_131_in_1, msg_to_bit_it_6_vnu_131_in_2, msg_to_bit_it_6_vnu_132_in_0, msg_to_bit_it_6_vnu_132_in_1, msg_to_bit_it_6_vnu_132_in_2, msg_to_bit_it_6_vnu_133_in_0, msg_to_bit_it_6_vnu_133_in_1, msg_to_bit_it_6_vnu_133_in_2, msg_to_bit_it_6_vnu_134_in_0, msg_to_bit_it_6_vnu_134_in_1, msg_to_bit_it_6_vnu_134_in_2, msg_to_bit_it_6_vnu_135_in_0, msg_to_bit_it_6_vnu_135_in_1, msg_to_bit_it_6_vnu_135_in_2, msg_to_bit_it_6_vnu_136_in_0, msg_to_bit_it_6_vnu_136_in_1, msg_to_bit_it_6_vnu_136_in_2, msg_to_bit_it_6_vnu_137_in_0, msg_to_bit_it_6_vnu_137_in_1, msg_to_bit_it_6_vnu_137_in_2, msg_to_bit_it_6_vnu_138_in_0, msg_to_bit_it_6_vnu_138_in_1, msg_to_bit_it_6_vnu_138_in_2, msg_to_bit_it_6_vnu_139_in_0, msg_to_bit_it_6_vnu_139_in_1, msg_to_bit_it_6_vnu_139_in_2, msg_to_bit_it_6_vnu_140_in_0, msg_to_bit_it_6_vnu_140_in_1, msg_to_bit_it_6_vnu_140_in_2, msg_to_bit_it_6_vnu_141_in_0, msg_to_bit_it_6_vnu_141_in_1, msg_to_bit_it_6_vnu_141_in_2, msg_to_bit_it_6_vnu_142_in_0, msg_to_bit_it_6_vnu_142_in_1, msg_to_bit_it_6_vnu_142_in_2, msg_to_bit_it_6_vnu_143_in_0, msg_to_bit_it_6_vnu_143_in_1, msg_to_bit_it_6_vnu_143_in_2, msg_to_bit_it_6_vnu_144_in_0, msg_to_bit_it_6_vnu_144_in_1, msg_to_bit_it_6_vnu_144_in_2, msg_to_bit_it_6_vnu_145_in_0, msg_to_bit_it_6_vnu_145_in_1, msg_to_bit_it_6_vnu_145_in_2, msg_to_bit_it_6_vnu_146_in_0, msg_to_bit_it_6_vnu_146_in_1, msg_to_bit_it_6_vnu_146_in_2, msg_to_bit_it_6_vnu_147_in_0, msg_to_bit_it_6_vnu_147_in_1, msg_to_bit_it_6_vnu_147_in_2, msg_to_bit_it_6_vnu_148_in_0, msg_to_bit_it_6_vnu_148_in_1, msg_to_bit_it_6_vnu_148_in_2, msg_to_bit_it_6_vnu_149_in_0, msg_to_bit_it_6_vnu_149_in_1, msg_to_bit_it_6_vnu_149_in_2, msg_to_bit_it_6_vnu_150_in_0, msg_to_bit_it_6_vnu_150_in_1, msg_to_bit_it_6_vnu_150_in_2, msg_to_bit_it_6_vnu_151_in_0, msg_to_bit_it_6_vnu_151_in_1, msg_to_bit_it_6_vnu_151_in_2, msg_to_bit_it_6_vnu_152_in_0, msg_to_bit_it_6_vnu_152_in_1, msg_to_bit_it_6_vnu_152_in_2, msg_to_bit_it_6_vnu_153_in_0, msg_to_bit_it_6_vnu_153_in_1, msg_to_bit_it_6_vnu_153_in_2, msg_to_bit_it_6_vnu_154_in_0, msg_to_bit_it_6_vnu_154_in_1, msg_to_bit_it_6_vnu_154_in_2, msg_to_bit_it_6_vnu_155_in_0, msg_to_bit_it_6_vnu_155_in_1, msg_to_bit_it_6_vnu_155_in_2, msg_to_bit_it_6_vnu_156_in_0, msg_to_bit_it_6_vnu_156_in_1, msg_to_bit_it_6_vnu_156_in_2, msg_to_bit_it_6_vnu_157_in_0, msg_to_bit_it_6_vnu_157_in_1, msg_to_bit_it_6_vnu_157_in_2, msg_to_bit_it_6_vnu_158_in_0, msg_to_bit_it_6_vnu_158_in_1, msg_to_bit_it_6_vnu_158_in_2, msg_to_bit_it_6_vnu_159_in_0, msg_to_bit_it_6_vnu_159_in_1, msg_to_bit_it_6_vnu_159_in_2, msg_to_bit_it_6_vnu_160_in_0, msg_to_bit_it_6_vnu_160_in_1, msg_to_bit_it_6_vnu_160_in_2, msg_to_bit_it_6_vnu_161_in_0, msg_to_bit_it_6_vnu_161_in_1, msg_to_bit_it_6_vnu_161_in_2, msg_to_bit_it_6_vnu_162_in_0, msg_to_bit_it_6_vnu_162_in_1, msg_to_bit_it_6_vnu_162_in_2, msg_to_bit_it_6_vnu_163_in_0, msg_to_bit_it_6_vnu_163_in_1, msg_to_bit_it_6_vnu_163_in_2, msg_to_bit_it_6_vnu_164_in_0, msg_to_bit_it_6_vnu_164_in_1, msg_to_bit_it_6_vnu_164_in_2, msg_to_bit_it_6_vnu_165_in_0, msg_to_bit_it_6_vnu_165_in_1, msg_to_bit_it_6_vnu_165_in_2, msg_to_bit_it_6_vnu_166_in_0, msg_to_bit_it_6_vnu_166_in_1, msg_to_bit_it_6_vnu_166_in_2, msg_to_bit_it_6_vnu_167_in_0, msg_to_bit_it_6_vnu_167_in_1, msg_to_bit_it_6_vnu_167_in_2, msg_to_bit_it_6_vnu_168_in_0, msg_to_bit_it_6_vnu_168_in_1, msg_to_bit_it_6_vnu_168_in_2, msg_to_bit_it_6_vnu_169_in_0, msg_to_bit_it_6_vnu_169_in_1, msg_to_bit_it_6_vnu_169_in_2, msg_to_bit_it_6_vnu_170_in_0, msg_to_bit_it_6_vnu_170_in_1, msg_to_bit_it_6_vnu_170_in_2, msg_to_bit_it_6_vnu_171_in_0, msg_to_bit_it_6_vnu_171_in_1, msg_to_bit_it_6_vnu_171_in_2, msg_to_bit_it_6_vnu_172_in_0, msg_to_bit_it_6_vnu_172_in_1, msg_to_bit_it_6_vnu_172_in_2, msg_to_bit_it_6_vnu_173_in_0, msg_to_bit_it_6_vnu_173_in_1, msg_to_bit_it_6_vnu_173_in_2, msg_to_bit_it_6_vnu_174_in_0, msg_to_bit_it_6_vnu_174_in_1, msg_to_bit_it_6_vnu_174_in_2, msg_to_bit_it_6_vnu_175_in_0, msg_to_bit_it_6_vnu_175_in_1, msg_to_bit_it_6_vnu_175_in_2, msg_to_bit_it_6_vnu_176_in_0, msg_to_bit_it_6_vnu_176_in_1, msg_to_bit_it_6_vnu_176_in_2, msg_to_bit_it_6_vnu_177_in_0, msg_to_bit_it_6_vnu_177_in_1, msg_to_bit_it_6_vnu_177_in_2, msg_to_bit_it_6_vnu_178_in_0, msg_to_bit_it_6_vnu_178_in_1, msg_to_bit_it_6_vnu_178_in_2, msg_to_bit_it_6_vnu_179_in_0, msg_to_bit_it_6_vnu_179_in_1, msg_to_bit_it_6_vnu_179_in_2, msg_to_bit_it_6_vnu_180_in_0, msg_to_bit_it_6_vnu_180_in_1, msg_to_bit_it_6_vnu_180_in_2, msg_to_bit_it_6_vnu_181_in_0, msg_to_bit_it_6_vnu_181_in_1, msg_to_bit_it_6_vnu_181_in_2, msg_to_bit_it_6_vnu_182_in_0, msg_to_bit_it_6_vnu_182_in_1, msg_to_bit_it_6_vnu_182_in_2, msg_to_bit_it_6_vnu_183_in_0, msg_to_bit_it_6_vnu_183_in_1, msg_to_bit_it_6_vnu_183_in_2, msg_to_bit_it_6_vnu_184_in_0, msg_to_bit_it_6_vnu_184_in_1, msg_to_bit_it_6_vnu_184_in_2, msg_to_bit_it_6_vnu_185_in_0, msg_to_bit_it_6_vnu_185_in_1, msg_to_bit_it_6_vnu_185_in_2, msg_to_bit_it_6_vnu_186_in_0, msg_to_bit_it_6_vnu_186_in_1, msg_to_bit_it_6_vnu_186_in_2, msg_to_bit_it_6_vnu_187_in_0, msg_to_bit_it_6_vnu_187_in_1, msg_to_bit_it_6_vnu_187_in_2, msg_to_bit_it_6_vnu_188_in_0, msg_to_bit_it_6_vnu_188_in_1, msg_to_bit_it_6_vnu_188_in_2, msg_to_bit_it_6_vnu_189_in_0, msg_to_bit_it_6_vnu_189_in_1, msg_to_bit_it_6_vnu_189_in_2, msg_to_bit_it_6_vnu_190_in_0, msg_to_bit_it_6_vnu_190_in_1, msg_to_bit_it_6_vnu_190_in_2, msg_to_bit_it_6_vnu_191_in_0, msg_to_bit_it_6_vnu_191_in_1, msg_to_bit_it_6_vnu_191_in_2, msg_to_bit_it_6_vnu_192_in_0, msg_to_bit_it_6_vnu_192_in_1, msg_to_bit_it_6_vnu_192_in_2, msg_to_bit_it_6_vnu_193_in_0, msg_to_bit_it_6_vnu_193_in_1, msg_to_bit_it_6_vnu_193_in_2, msg_to_bit_it_6_vnu_194_in_0, msg_to_bit_it_6_vnu_194_in_1, msg_to_bit_it_6_vnu_194_in_2, msg_to_bit_it_6_vnu_195_in_0, msg_to_bit_it_6_vnu_195_in_1, msg_to_bit_it_6_vnu_195_in_2, msg_to_bit_it_6_vnu_196_in_0, msg_to_bit_it_6_vnu_196_in_1, msg_to_bit_it_6_vnu_196_in_2, msg_to_bit_it_6_vnu_197_in_0, msg_to_bit_it_6_vnu_197_in_1, msg_to_bit_it_6_vnu_197_in_2, msg_to_bit_it_7_vnu_0_in_0, msg_to_bit_it_7_vnu_0_in_1, msg_to_bit_it_7_vnu_0_in_2, msg_to_bit_it_7_vnu_1_in_0, msg_to_bit_it_7_vnu_1_in_1, msg_to_bit_it_7_vnu_1_in_2, msg_to_bit_it_7_vnu_2_in_0, msg_to_bit_it_7_vnu_2_in_1, msg_to_bit_it_7_vnu_2_in_2, msg_to_bit_it_7_vnu_3_in_0, msg_to_bit_it_7_vnu_3_in_1, msg_to_bit_it_7_vnu_3_in_2, msg_to_bit_it_7_vnu_4_in_0, msg_to_bit_it_7_vnu_4_in_1, msg_to_bit_it_7_vnu_4_in_2, msg_to_bit_it_7_vnu_5_in_0, msg_to_bit_it_7_vnu_5_in_1, msg_to_bit_it_7_vnu_5_in_2, msg_to_bit_it_7_vnu_6_in_0, msg_to_bit_it_7_vnu_6_in_1, msg_to_bit_it_7_vnu_6_in_2, msg_to_bit_it_7_vnu_7_in_0, msg_to_bit_it_7_vnu_7_in_1, msg_to_bit_it_7_vnu_7_in_2, msg_to_bit_it_7_vnu_8_in_0, msg_to_bit_it_7_vnu_8_in_1, msg_to_bit_it_7_vnu_8_in_2, msg_to_bit_it_7_vnu_9_in_0, msg_to_bit_it_7_vnu_9_in_1, msg_to_bit_it_7_vnu_9_in_2, msg_to_bit_it_7_vnu_10_in_0, msg_to_bit_it_7_vnu_10_in_1, msg_to_bit_it_7_vnu_10_in_2, msg_to_bit_it_7_vnu_11_in_0, msg_to_bit_it_7_vnu_11_in_1, msg_to_bit_it_7_vnu_11_in_2, msg_to_bit_it_7_vnu_12_in_0, msg_to_bit_it_7_vnu_12_in_1, msg_to_bit_it_7_vnu_12_in_2, msg_to_bit_it_7_vnu_13_in_0, msg_to_bit_it_7_vnu_13_in_1, msg_to_bit_it_7_vnu_13_in_2, msg_to_bit_it_7_vnu_14_in_0, msg_to_bit_it_7_vnu_14_in_1, msg_to_bit_it_7_vnu_14_in_2, msg_to_bit_it_7_vnu_15_in_0, msg_to_bit_it_7_vnu_15_in_1, msg_to_bit_it_7_vnu_15_in_2, msg_to_bit_it_7_vnu_16_in_0, msg_to_bit_it_7_vnu_16_in_1, msg_to_bit_it_7_vnu_16_in_2, msg_to_bit_it_7_vnu_17_in_0, msg_to_bit_it_7_vnu_17_in_1, msg_to_bit_it_7_vnu_17_in_2, msg_to_bit_it_7_vnu_18_in_0, msg_to_bit_it_7_vnu_18_in_1, msg_to_bit_it_7_vnu_18_in_2, msg_to_bit_it_7_vnu_19_in_0, msg_to_bit_it_7_vnu_19_in_1, msg_to_bit_it_7_vnu_19_in_2, msg_to_bit_it_7_vnu_20_in_0, msg_to_bit_it_7_vnu_20_in_1, msg_to_bit_it_7_vnu_20_in_2, msg_to_bit_it_7_vnu_21_in_0, msg_to_bit_it_7_vnu_21_in_1, msg_to_bit_it_7_vnu_21_in_2, msg_to_bit_it_7_vnu_22_in_0, msg_to_bit_it_7_vnu_22_in_1, msg_to_bit_it_7_vnu_22_in_2, msg_to_bit_it_7_vnu_23_in_0, msg_to_bit_it_7_vnu_23_in_1, msg_to_bit_it_7_vnu_23_in_2, msg_to_bit_it_7_vnu_24_in_0, msg_to_bit_it_7_vnu_24_in_1, msg_to_bit_it_7_vnu_24_in_2, msg_to_bit_it_7_vnu_25_in_0, msg_to_bit_it_7_vnu_25_in_1, msg_to_bit_it_7_vnu_25_in_2, msg_to_bit_it_7_vnu_26_in_0, msg_to_bit_it_7_vnu_26_in_1, msg_to_bit_it_7_vnu_26_in_2, msg_to_bit_it_7_vnu_27_in_0, msg_to_bit_it_7_vnu_27_in_1, msg_to_bit_it_7_vnu_27_in_2, msg_to_bit_it_7_vnu_28_in_0, msg_to_bit_it_7_vnu_28_in_1, msg_to_bit_it_7_vnu_28_in_2, msg_to_bit_it_7_vnu_29_in_0, msg_to_bit_it_7_vnu_29_in_1, msg_to_bit_it_7_vnu_29_in_2, msg_to_bit_it_7_vnu_30_in_0, msg_to_bit_it_7_vnu_30_in_1, msg_to_bit_it_7_vnu_30_in_2, msg_to_bit_it_7_vnu_31_in_0, msg_to_bit_it_7_vnu_31_in_1, msg_to_bit_it_7_vnu_31_in_2, msg_to_bit_it_7_vnu_32_in_0, msg_to_bit_it_7_vnu_32_in_1, msg_to_bit_it_7_vnu_32_in_2, msg_to_bit_it_7_vnu_33_in_0, msg_to_bit_it_7_vnu_33_in_1, msg_to_bit_it_7_vnu_33_in_2, msg_to_bit_it_7_vnu_34_in_0, msg_to_bit_it_7_vnu_34_in_1, msg_to_bit_it_7_vnu_34_in_2, msg_to_bit_it_7_vnu_35_in_0, msg_to_bit_it_7_vnu_35_in_1, msg_to_bit_it_7_vnu_35_in_2, msg_to_bit_it_7_vnu_36_in_0, msg_to_bit_it_7_vnu_36_in_1, msg_to_bit_it_7_vnu_36_in_2, msg_to_bit_it_7_vnu_37_in_0, msg_to_bit_it_7_vnu_37_in_1, msg_to_bit_it_7_vnu_37_in_2, msg_to_bit_it_7_vnu_38_in_0, msg_to_bit_it_7_vnu_38_in_1, msg_to_bit_it_7_vnu_38_in_2, msg_to_bit_it_7_vnu_39_in_0, msg_to_bit_it_7_vnu_39_in_1, msg_to_bit_it_7_vnu_39_in_2, msg_to_bit_it_7_vnu_40_in_0, msg_to_bit_it_7_vnu_40_in_1, msg_to_bit_it_7_vnu_40_in_2, msg_to_bit_it_7_vnu_41_in_0, msg_to_bit_it_7_vnu_41_in_1, msg_to_bit_it_7_vnu_41_in_2, msg_to_bit_it_7_vnu_42_in_0, msg_to_bit_it_7_vnu_42_in_1, msg_to_bit_it_7_vnu_42_in_2, msg_to_bit_it_7_vnu_43_in_0, msg_to_bit_it_7_vnu_43_in_1, msg_to_bit_it_7_vnu_43_in_2, msg_to_bit_it_7_vnu_44_in_0, msg_to_bit_it_7_vnu_44_in_1, msg_to_bit_it_7_vnu_44_in_2, msg_to_bit_it_7_vnu_45_in_0, msg_to_bit_it_7_vnu_45_in_1, msg_to_bit_it_7_vnu_45_in_2, msg_to_bit_it_7_vnu_46_in_0, msg_to_bit_it_7_vnu_46_in_1, msg_to_bit_it_7_vnu_46_in_2, msg_to_bit_it_7_vnu_47_in_0, msg_to_bit_it_7_vnu_47_in_1, msg_to_bit_it_7_vnu_47_in_2, msg_to_bit_it_7_vnu_48_in_0, msg_to_bit_it_7_vnu_48_in_1, msg_to_bit_it_7_vnu_48_in_2, msg_to_bit_it_7_vnu_49_in_0, msg_to_bit_it_7_vnu_49_in_1, msg_to_bit_it_7_vnu_49_in_2, msg_to_bit_it_7_vnu_50_in_0, msg_to_bit_it_7_vnu_50_in_1, msg_to_bit_it_7_vnu_50_in_2, msg_to_bit_it_7_vnu_51_in_0, msg_to_bit_it_7_vnu_51_in_1, msg_to_bit_it_7_vnu_51_in_2, msg_to_bit_it_7_vnu_52_in_0, msg_to_bit_it_7_vnu_52_in_1, msg_to_bit_it_7_vnu_52_in_2, msg_to_bit_it_7_vnu_53_in_0, msg_to_bit_it_7_vnu_53_in_1, msg_to_bit_it_7_vnu_53_in_2, msg_to_bit_it_7_vnu_54_in_0, msg_to_bit_it_7_vnu_54_in_1, msg_to_bit_it_7_vnu_54_in_2, msg_to_bit_it_7_vnu_55_in_0, msg_to_bit_it_7_vnu_55_in_1, msg_to_bit_it_7_vnu_55_in_2, msg_to_bit_it_7_vnu_56_in_0, msg_to_bit_it_7_vnu_56_in_1, msg_to_bit_it_7_vnu_56_in_2, msg_to_bit_it_7_vnu_57_in_0, msg_to_bit_it_7_vnu_57_in_1, msg_to_bit_it_7_vnu_57_in_2, msg_to_bit_it_7_vnu_58_in_0, msg_to_bit_it_7_vnu_58_in_1, msg_to_bit_it_7_vnu_58_in_2, msg_to_bit_it_7_vnu_59_in_0, msg_to_bit_it_7_vnu_59_in_1, msg_to_bit_it_7_vnu_59_in_2, msg_to_bit_it_7_vnu_60_in_0, msg_to_bit_it_7_vnu_60_in_1, msg_to_bit_it_7_vnu_60_in_2, msg_to_bit_it_7_vnu_61_in_0, msg_to_bit_it_7_vnu_61_in_1, msg_to_bit_it_7_vnu_61_in_2, msg_to_bit_it_7_vnu_62_in_0, msg_to_bit_it_7_vnu_62_in_1, msg_to_bit_it_7_vnu_62_in_2, msg_to_bit_it_7_vnu_63_in_0, msg_to_bit_it_7_vnu_63_in_1, msg_to_bit_it_7_vnu_63_in_2, msg_to_bit_it_7_vnu_64_in_0, msg_to_bit_it_7_vnu_64_in_1, msg_to_bit_it_7_vnu_64_in_2, msg_to_bit_it_7_vnu_65_in_0, msg_to_bit_it_7_vnu_65_in_1, msg_to_bit_it_7_vnu_65_in_2, msg_to_bit_it_7_vnu_66_in_0, msg_to_bit_it_7_vnu_66_in_1, msg_to_bit_it_7_vnu_66_in_2, msg_to_bit_it_7_vnu_67_in_0, msg_to_bit_it_7_vnu_67_in_1, msg_to_bit_it_7_vnu_67_in_2, msg_to_bit_it_7_vnu_68_in_0, msg_to_bit_it_7_vnu_68_in_1, msg_to_bit_it_7_vnu_68_in_2, msg_to_bit_it_7_vnu_69_in_0, msg_to_bit_it_7_vnu_69_in_1, msg_to_bit_it_7_vnu_69_in_2, msg_to_bit_it_7_vnu_70_in_0, msg_to_bit_it_7_vnu_70_in_1, msg_to_bit_it_7_vnu_70_in_2, msg_to_bit_it_7_vnu_71_in_0, msg_to_bit_it_7_vnu_71_in_1, msg_to_bit_it_7_vnu_71_in_2, msg_to_bit_it_7_vnu_72_in_0, msg_to_bit_it_7_vnu_72_in_1, msg_to_bit_it_7_vnu_72_in_2, msg_to_bit_it_7_vnu_73_in_0, msg_to_bit_it_7_vnu_73_in_1, msg_to_bit_it_7_vnu_73_in_2, msg_to_bit_it_7_vnu_74_in_0, msg_to_bit_it_7_vnu_74_in_1, msg_to_bit_it_7_vnu_74_in_2, msg_to_bit_it_7_vnu_75_in_0, msg_to_bit_it_7_vnu_75_in_1, msg_to_bit_it_7_vnu_75_in_2, msg_to_bit_it_7_vnu_76_in_0, msg_to_bit_it_7_vnu_76_in_1, msg_to_bit_it_7_vnu_76_in_2, msg_to_bit_it_7_vnu_77_in_0, msg_to_bit_it_7_vnu_77_in_1, msg_to_bit_it_7_vnu_77_in_2, msg_to_bit_it_7_vnu_78_in_0, msg_to_bit_it_7_vnu_78_in_1, msg_to_bit_it_7_vnu_78_in_2, msg_to_bit_it_7_vnu_79_in_0, msg_to_bit_it_7_vnu_79_in_1, msg_to_bit_it_7_vnu_79_in_2, msg_to_bit_it_7_vnu_80_in_0, msg_to_bit_it_7_vnu_80_in_1, msg_to_bit_it_7_vnu_80_in_2, msg_to_bit_it_7_vnu_81_in_0, msg_to_bit_it_7_vnu_81_in_1, msg_to_bit_it_7_vnu_81_in_2, msg_to_bit_it_7_vnu_82_in_0, msg_to_bit_it_7_vnu_82_in_1, msg_to_bit_it_7_vnu_82_in_2, msg_to_bit_it_7_vnu_83_in_0, msg_to_bit_it_7_vnu_83_in_1, msg_to_bit_it_7_vnu_83_in_2, msg_to_bit_it_7_vnu_84_in_0, msg_to_bit_it_7_vnu_84_in_1, msg_to_bit_it_7_vnu_84_in_2, msg_to_bit_it_7_vnu_85_in_0, msg_to_bit_it_7_vnu_85_in_1, msg_to_bit_it_7_vnu_85_in_2, msg_to_bit_it_7_vnu_86_in_0, msg_to_bit_it_7_vnu_86_in_1, msg_to_bit_it_7_vnu_86_in_2, msg_to_bit_it_7_vnu_87_in_0, msg_to_bit_it_7_vnu_87_in_1, msg_to_bit_it_7_vnu_87_in_2, msg_to_bit_it_7_vnu_88_in_0, msg_to_bit_it_7_vnu_88_in_1, msg_to_bit_it_7_vnu_88_in_2, msg_to_bit_it_7_vnu_89_in_0, msg_to_bit_it_7_vnu_89_in_1, msg_to_bit_it_7_vnu_89_in_2, msg_to_bit_it_7_vnu_90_in_0, msg_to_bit_it_7_vnu_90_in_1, msg_to_bit_it_7_vnu_90_in_2, msg_to_bit_it_7_vnu_91_in_0, msg_to_bit_it_7_vnu_91_in_1, msg_to_bit_it_7_vnu_91_in_2, msg_to_bit_it_7_vnu_92_in_0, msg_to_bit_it_7_vnu_92_in_1, msg_to_bit_it_7_vnu_92_in_2, msg_to_bit_it_7_vnu_93_in_0, msg_to_bit_it_7_vnu_93_in_1, msg_to_bit_it_7_vnu_93_in_2, msg_to_bit_it_7_vnu_94_in_0, msg_to_bit_it_7_vnu_94_in_1, msg_to_bit_it_7_vnu_94_in_2, msg_to_bit_it_7_vnu_95_in_0, msg_to_bit_it_7_vnu_95_in_1, msg_to_bit_it_7_vnu_95_in_2, msg_to_bit_it_7_vnu_96_in_0, msg_to_bit_it_7_vnu_96_in_1, msg_to_bit_it_7_vnu_96_in_2, msg_to_bit_it_7_vnu_97_in_0, msg_to_bit_it_7_vnu_97_in_1, msg_to_bit_it_7_vnu_97_in_2, msg_to_bit_it_7_vnu_98_in_0, msg_to_bit_it_7_vnu_98_in_1, msg_to_bit_it_7_vnu_98_in_2, msg_to_bit_it_7_vnu_99_in_0, msg_to_bit_it_7_vnu_99_in_1, msg_to_bit_it_7_vnu_99_in_2, msg_to_bit_it_7_vnu_100_in_0, msg_to_bit_it_7_vnu_100_in_1, msg_to_bit_it_7_vnu_100_in_2, msg_to_bit_it_7_vnu_101_in_0, msg_to_bit_it_7_vnu_101_in_1, msg_to_bit_it_7_vnu_101_in_2, msg_to_bit_it_7_vnu_102_in_0, msg_to_bit_it_7_vnu_102_in_1, msg_to_bit_it_7_vnu_102_in_2, msg_to_bit_it_7_vnu_103_in_0, msg_to_bit_it_7_vnu_103_in_1, msg_to_bit_it_7_vnu_103_in_2, msg_to_bit_it_7_vnu_104_in_0, msg_to_bit_it_7_vnu_104_in_1, msg_to_bit_it_7_vnu_104_in_2, msg_to_bit_it_7_vnu_105_in_0, msg_to_bit_it_7_vnu_105_in_1, msg_to_bit_it_7_vnu_105_in_2, msg_to_bit_it_7_vnu_106_in_0, msg_to_bit_it_7_vnu_106_in_1, msg_to_bit_it_7_vnu_106_in_2, msg_to_bit_it_7_vnu_107_in_0, msg_to_bit_it_7_vnu_107_in_1, msg_to_bit_it_7_vnu_107_in_2, msg_to_bit_it_7_vnu_108_in_0, msg_to_bit_it_7_vnu_108_in_1, msg_to_bit_it_7_vnu_108_in_2, msg_to_bit_it_7_vnu_109_in_0, msg_to_bit_it_7_vnu_109_in_1, msg_to_bit_it_7_vnu_109_in_2, msg_to_bit_it_7_vnu_110_in_0, msg_to_bit_it_7_vnu_110_in_1, msg_to_bit_it_7_vnu_110_in_2, msg_to_bit_it_7_vnu_111_in_0, msg_to_bit_it_7_vnu_111_in_1, msg_to_bit_it_7_vnu_111_in_2, msg_to_bit_it_7_vnu_112_in_0, msg_to_bit_it_7_vnu_112_in_1, msg_to_bit_it_7_vnu_112_in_2, msg_to_bit_it_7_vnu_113_in_0, msg_to_bit_it_7_vnu_113_in_1, msg_to_bit_it_7_vnu_113_in_2, msg_to_bit_it_7_vnu_114_in_0, msg_to_bit_it_7_vnu_114_in_1, msg_to_bit_it_7_vnu_114_in_2, msg_to_bit_it_7_vnu_115_in_0, msg_to_bit_it_7_vnu_115_in_1, msg_to_bit_it_7_vnu_115_in_2, msg_to_bit_it_7_vnu_116_in_0, msg_to_bit_it_7_vnu_116_in_1, msg_to_bit_it_7_vnu_116_in_2, msg_to_bit_it_7_vnu_117_in_0, msg_to_bit_it_7_vnu_117_in_1, msg_to_bit_it_7_vnu_117_in_2, msg_to_bit_it_7_vnu_118_in_0, msg_to_bit_it_7_vnu_118_in_1, msg_to_bit_it_7_vnu_118_in_2, msg_to_bit_it_7_vnu_119_in_0, msg_to_bit_it_7_vnu_119_in_1, msg_to_bit_it_7_vnu_119_in_2, msg_to_bit_it_7_vnu_120_in_0, msg_to_bit_it_7_vnu_120_in_1, msg_to_bit_it_7_vnu_120_in_2, msg_to_bit_it_7_vnu_121_in_0, msg_to_bit_it_7_vnu_121_in_1, msg_to_bit_it_7_vnu_121_in_2, msg_to_bit_it_7_vnu_122_in_0, msg_to_bit_it_7_vnu_122_in_1, msg_to_bit_it_7_vnu_122_in_2, msg_to_bit_it_7_vnu_123_in_0, msg_to_bit_it_7_vnu_123_in_1, msg_to_bit_it_7_vnu_123_in_2, msg_to_bit_it_7_vnu_124_in_0, msg_to_bit_it_7_vnu_124_in_1, msg_to_bit_it_7_vnu_124_in_2, msg_to_bit_it_7_vnu_125_in_0, msg_to_bit_it_7_vnu_125_in_1, msg_to_bit_it_7_vnu_125_in_2, msg_to_bit_it_7_vnu_126_in_0, msg_to_bit_it_7_vnu_126_in_1, msg_to_bit_it_7_vnu_126_in_2, msg_to_bit_it_7_vnu_127_in_0, msg_to_bit_it_7_vnu_127_in_1, msg_to_bit_it_7_vnu_127_in_2, msg_to_bit_it_7_vnu_128_in_0, msg_to_bit_it_7_vnu_128_in_1, msg_to_bit_it_7_vnu_128_in_2, msg_to_bit_it_7_vnu_129_in_0, msg_to_bit_it_7_vnu_129_in_1, msg_to_bit_it_7_vnu_129_in_2, msg_to_bit_it_7_vnu_130_in_0, msg_to_bit_it_7_vnu_130_in_1, msg_to_bit_it_7_vnu_130_in_2, msg_to_bit_it_7_vnu_131_in_0, msg_to_bit_it_7_vnu_131_in_1, msg_to_bit_it_7_vnu_131_in_2, msg_to_bit_it_7_vnu_132_in_0, msg_to_bit_it_7_vnu_132_in_1, msg_to_bit_it_7_vnu_132_in_2, msg_to_bit_it_7_vnu_133_in_0, msg_to_bit_it_7_vnu_133_in_1, msg_to_bit_it_7_vnu_133_in_2, msg_to_bit_it_7_vnu_134_in_0, msg_to_bit_it_7_vnu_134_in_1, msg_to_bit_it_7_vnu_134_in_2, msg_to_bit_it_7_vnu_135_in_0, msg_to_bit_it_7_vnu_135_in_1, msg_to_bit_it_7_vnu_135_in_2, msg_to_bit_it_7_vnu_136_in_0, msg_to_bit_it_7_vnu_136_in_1, msg_to_bit_it_7_vnu_136_in_2, msg_to_bit_it_7_vnu_137_in_0, msg_to_bit_it_7_vnu_137_in_1, msg_to_bit_it_7_vnu_137_in_2, msg_to_bit_it_7_vnu_138_in_0, msg_to_bit_it_7_vnu_138_in_1, msg_to_bit_it_7_vnu_138_in_2, msg_to_bit_it_7_vnu_139_in_0, msg_to_bit_it_7_vnu_139_in_1, msg_to_bit_it_7_vnu_139_in_2, msg_to_bit_it_7_vnu_140_in_0, msg_to_bit_it_7_vnu_140_in_1, msg_to_bit_it_7_vnu_140_in_2, msg_to_bit_it_7_vnu_141_in_0, msg_to_bit_it_7_vnu_141_in_1, msg_to_bit_it_7_vnu_141_in_2, msg_to_bit_it_7_vnu_142_in_0, msg_to_bit_it_7_vnu_142_in_1, msg_to_bit_it_7_vnu_142_in_2, msg_to_bit_it_7_vnu_143_in_0, msg_to_bit_it_7_vnu_143_in_1, msg_to_bit_it_7_vnu_143_in_2, msg_to_bit_it_7_vnu_144_in_0, msg_to_bit_it_7_vnu_144_in_1, msg_to_bit_it_7_vnu_144_in_2, msg_to_bit_it_7_vnu_145_in_0, msg_to_bit_it_7_vnu_145_in_1, msg_to_bit_it_7_vnu_145_in_2, msg_to_bit_it_7_vnu_146_in_0, msg_to_bit_it_7_vnu_146_in_1, msg_to_bit_it_7_vnu_146_in_2, msg_to_bit_it_7_vnu_147_in_0, msg_to_bit_it_7_vnu_147_in_1, msg_to_bit_it_7_vnu_147_in_2, msg_to_bit_it_7_vnu_148_in_0, msg_to_bit_it_7_vnu_148_in_1, msg_to_bit_it_7_vnu_148_in_2, msg_to_bit_it_7_vnu_149_in_0, msg_to_bit_it_7_vnu_149_in_1, msg_to_bit_it_7_vnu_149_in_2, msg_to_bit_it_7_vnu_150_in_0, msg_to_bit_it_7_vnu_150_in_1, msg_to_bit_it_7_vnu_150_in_2, msg_to_bit_it_7_vnu_151_in_0, msg_to_bit_it_7_vnu_151_in_1, msg_to_bit_it_7_vnu_151_in_2, msg_to_bit_it_7_vnu_152_in_0, msg_to_bit_it_7_vnu_152_in_1, msg_to_bit_it_7_vnu_152_in_2, msg_to_bit_it_7_vnu_153_in_0, msg_to_bit_it_7_vnu_153_in_1, msg_to_bit_it_7_vnu_153_in_2, msg_to_bit_it_7_vnu_154_in_0, msg_to_bit_it_7_vnu_154_in_1, msg_to_bit_it_7_vnu_154_in_2, msg_to_bit_it_7_vnu_155_in_0, msg_to_bit_it_7_vnu_155_in_1, msg_to_bit_it_7_vnu_155_in_2, msg_to_bit_it_7_vnu_156_in_0, msg_to_bit_it_7_vnu_156_in_1, msg_to_bit_it_7_vnu_156_in_2, msg_to_bit_it_7_vnu_157_in_0, msg_to_bit_it_7_vnu_157_in_1, msg_to_bit_it_7_vnu_157_in_2, msg_to_bit_it_7_vnu_158_in_0, msg_to_bit_it_7_vnu_158_in_1, msg_to_bit_it_7_vnu_158_in_2, msg_to_bit_it_7_vnu_159_in_0, msg_to_bit_it_7_vnu_159_in_1, msg_to_bit_it_7_vnu_159_in_2, msg_to_bit_it_7_vnu_160_in_0, msg_to_bit_it_7_vnu_160_in_1, msg_to_bit_it_7_vnu_160_in_2, msg_to_bit_it_7_vnu_161_in_0, msg_to_bit_it_7_vnu_161_in_1, msg_to_bit_it_7_vnu_161_in_2, msg_to_bit_it_7_vnu_162_in_0, msg_to_bit_it_7_vnu_162_in_1, msg_to_bit_it_7_vnu_162_in_2, msg_to_bit_it_7_vnu_163_in_0, msg_to_bit_it_7_vnu_163_in_1, msg_to_bit_it_7_vnu_163_in_2, msg_to_bit_it_7_vnu_164_in_0, msg_to_bit_it_7_vnu_164_in_1, msg_to_bit_it_7_vnu_164_in_2, msg_to_bit_it_7_vnu_165_in_0, msg_to_bit_it_7_vnu_165_in_1, msg_to_bit_it_7_vnu_165_in_2, msg_to_bit_it_7_vnu_166_in_0, msg_to_bit_it_7_vnu_166_in_1, msg_to_bit_it_7_vnu_166_in_2, msg_to_bit_it_7_vnu_167_in_0, msg_to_bit_it_7_vnu_167_in_1, msg_to_bit_it_7_vnu_167_in_2, msg_to_bit_it_7_vnu_168_in_0, msg_to_bit_it_7_vnu_168_in_1, msg_to_bit_it_7_vnu_168_in_2, msg_to_bit_it_7_vnu_169_in_0, msg_to_bit_it_7_vnu_169_in_1, msg_to_bit_it_7_vnu_169_in_2, msg_to_bit_it_7_vnu_170_in_0, msg_to_bit_it_7_vnu_170_in_1, msg_to_bit_it_7_vnu_170_in_2, msg_to_bit_it_7_vnu_171_in_0, msg_to_bit_it_7_vnu_171_in_1, msg_to_bit_it_7_vnu_171_in_2, msg_to_bit_it_7_vnu_172_in_0, msg_to_bit_it_7_vnu_172_in_1, msg_to_bit_it_7_vnu_172_in_2, msg_to_bit_it_7_vnu_173_in_0, msg_to_bit_it_7_vnu_173_in_1, msg_to_bit_it_7_vnu_173_in_2, msg_to_bit_it_7_vnu_174_in_0, msg_to_bit_it_7_vnu_174_in_1, msg_to_bit_it_7_vnu_174_in_2, msg_to_bit_it_7_vnu_175_in_0, msg_to_bit_it_7_vnu_175_in_1, msg_to_bit_it_7_vnu_175_in_2, msg_to_bit_it_7_vnu_176_in_0, msg_to_bit_it_7_vnu_176_in_1, msg_to_bit_it_7_vnu_176_in_2, msg_to_bit_it_7_vnu_177_in_0, msg_to_bit_it_7_vnu_177_in_1, msg_to_bit_it_7_vnu_177_in_2, msg_to_bit_it_7_vnu_178_in_0, msg_to_bit_it_7_vnu_178_in_1, msg_to_bit_it_7_vnu_178_in_2, msg_to_bit_it_7_vnu_179_in_0, msg_to_bit_it_7_vnu_179_in_1, msg_to_bit_it_7_vnu_179_in_2, msg_to_bit_it_7_vnu_180_in_0, msg_to_bit_it_7_vnu_180_in_1, msg_to_bit_it_7_vnu_180_in_2, msg_to_bit_it_7_vnu_181_in_0, msg_to_bit_it_7_vnu_181_in_1, msg_to_bit_it_7_vnu_181_in_2, msg_to_bit_it_7_vnu_182_in_0, msg_to_bit_it_7_vnu_182_in_1, msg_to_bit_it_7_vnu_182_in_2, msg_to_bit_it_7_vnu_183_in_0, msg_to_bit_it_7_vnu_183_in_1, msg_to_bit_it_7_vnu_183_in_2, msg_to_bit_it_7_vnu_184_in_0, msg_to_bit_it_7_vnu_184_in_1, msg_to_bit_it_7_vnu_184_in_2, msg_to_bit_it_7_vnu_185_in_0, msg_to_bit_it_7_vnu_185_in_1, msg_to_bit_it_7_vnu_185_in_2, msg_to_bit_it_7_vnu_186_in_0, msg_to_bit_it_7_vnu_186_in_1, msg_to_bit_it_7_vnu_186_in_2, msg_to_bit_it_7_vnu_187_in_0, msg_to_bit_it_7_vnu_187_in_1, msg_to_bit_it_7_vnu_187_in_2, msg_to_bit_it_7_vnu_188_in_0, msg_to_bit_it_7_vnu_188_in_1, msg_to_bit_it_7_vnu_188_in_2, msg_to_bit_it_7_vnu_189_in_0, msg_to_bit_it_7_vnu_189_in_1, msg_to_bit_it_7_vnu_189_in_2, msg_to_bit_it_7_vnu_190_in_0, msg_to_bit_it_7_vnu_190_in_1, msg_to_bit_it_7_vnu_190_in_2, msg_to_bit_it_7_vnu_191_in_0, msg_to_bit_it_7_vnu_191_in_1, msg_to_bit_it_7_vnu_191_in_2, msg_to_bit_it_7_vnu_192_in_0, msg_to_bit_it_7_vnu_192_in_1, msg_to_bit_it_7_vnu_192_in_2, msg_to_bit_it_7_vnu_193_in_0, msg_to_bit_it_7_vnu_193_in_1, msg_to_bit_it_7_vnu_193_in_2, msg_to_bit_it_7_vnu_194_in_0, msg_to_bit_it_7_vnu_194_in_1, msg_to_bit_it_7_vnu_194_in_2, msg_to_bit_it_7_vnu_195_in_0, msg_to_bit_it_7_vnu_195_in_1, msg_to_bit_it_7_vnu_195_in_2, msg_to_bit_it_7_vnu_196_in_0, msg_to_bit_it_7_vnu_196_in_1, msg_to_bit_it_7_vnu_196_in_2, msg_to_bit_it_7_vnu_197_in_0, msg_to_bit_it_7_vnu_197_in_1, msg_to_bit_it_7_vnu_197_in_2, msg_to_bit_it_8_vnu_0_in_0, msg_to_bit_it_8_vnu_0_in_1, msg_to_bit_it_8_vnu_0_in_2, msg_to_bit_it_8_vnu_1_in_0, msg_to_bit_it_8_vnu_1_in_1, msg_to_bit_it_8_vnu_1_in_2, msg_to_bit_it_8_vnu_2_in_0, msg_to_bit_it_8_vnu_2_in_1, msg_to_bit_it_8_vnu_2_in_2, msg_to_bit_it_8_vnu_3_in_0, msg_to_bit_it_8_vnu_3_in_1, msg_to_bit_it_8_vnu_3_in_2, msg_to_bit_it_8_vnu_4_in_0, msg_to_bit_it_8_vnu_4_in_1, msg_to_bit_it_8_vnu_4_in_2, msg_to_bit_it_8_vnu_5_in_0, msg_to_bit_it_8_vnu_5_in_1, msg_to_bit_it_8_vnu_5_in_2, msg_to_bit_it_8_vnu_6_in_0, msg_to_bit_it_8_vnu_6_in_1, msg_to_bit_it_8_vnu_6_in_2, msg_to_bit_it_8_vnu_7_in_0, msg_to_bit_it_8_vnu_7_in_1, msg_to_bit_it_8_vnu_7_in_2, msg_to_bit_it_8_vnu_8_in_0, msg_to_bit_it_8_vnu_8_in_1, msg_to_bit_it_8_vnu_8_in_2, msg_to_bit_it_8_vnu_9_in_0, msg_to_bit_it_8_vnu_9_in_1, msg_to_bit_it_8_vnu_9_in_2, msg_to_bit_it_8_vnu_10_in_0, msg_to_bit_it_8_vnu_10_in_1, msg_to_bit_it_8_vnu_10_in_2, msg_to_bit_it_8_vnu_11_in_0, msg_to_bit_it_8_vnu_11_in_1, msg_to_bit_it_8_vnu_11_in_2, msg_to_bit_it_8_vnu_12_in_0, msg_to_bit_it_8_vnu_12_in_1, msg_to_bit_it_8_vnu_12_in_2, msg_to_bit_it_8_vnu_13_in_0, msg_to_bit_it_8_vnu_13_in_1, msg_to_bit_it_8_vnu_13_in_2, msg_to_bit_it_8_vnu_14_in_0, msg_to_bit_it_8_vnu_14_in_1, msg_to_bit_it_8_vnu_14_in_2, msg_to_bit_it_8_vnu_15_in_0, msg_to_bit_it_8_vnu_15_in_1, msg_to_bit_it_8_vnu_15_in_2, msg_to_bit_it_8_vnu_16_in_0, msg_to_bit_it_8_vnu_16_in_1, msg_to_bit_it_8_vnu_16_in_2, msg_to_bit_it_8_vnu_17_in_0, msg_to_bit_it_8_vnu_17_in_1, msg_to_bit_it_8_vnu_17_in_2, msg_to_bit_it_8_vnu_18_in_0, msg_to_bit_it_8_vnu_18_in_1, msg_to_bit_it_8_vnu_18_in_2, msg_to_bit_it_8_vnu_19_in_0, msg_to_bit_it_8_vnu_19_in_1, msg_to_bit_it_8_vnu_19_in_2, msg_to_bit_it_8_vnu_20_in_0, msg_to_bit_it_8_vnu_20_in_1, msg_to_bit_it_8_vnu_20_in_2, msg_to_bit_it_8_vnu_21_in_0, msg_to_bit_it_8_vnu_21_in_1, msg_to_bit_it_8_vnu_21_in_2, msg_to_bit_it_8_vnu_22_in_0, msg_to_bit_it_8_vnu_22_in_1, msg_to_bit_it_8_vnu_22_in_2, msg_to_bit_it_8_vnu_23_in_0, msg_to_bit_it_8_vnu_23_in_1, msg_to_bit_it_8_vnu_23_in_2, msg_to_bit_it_8_vnu_24_in_0, msg_to_bit_it_8_vnu_24_in_1, msg_to_bit_it_8_vnu_24_in_2, msg_to_bit_it_8_vnu_25_in_0, msg_to_bit_it_8_vnu_25_in_1, msg_to_bit_it_8_vnu_25_in_2, msg_to_bit_it_8_vnu_26_in_0, msg_to_bit_it_8_vnu_26_in_1, msg_to_bit_it_8_vnu_26_in_2, msg_to_bit_it_8_vnu_27_in_0, msg_to_bit_it_8_vnu_27_in_1, msg_to_bit_it_8_vnu_27_in_2, msg_to_bit_it_8_vnu_28_in_0, msg_to_bit_it_8_vnu_28_in_1, msg_to_bit_it_8_vnu_28_in_2, msg_to_bit_it_8_vnu_29_in_0, msg_to_bit_it_8_vnu_29_in_1, msg_to_bit_it_8_vnu_29_in_2, msg_to_bit_it_8_vnu_30_in_0, msg_to_bit_it_8_vnu_30_in_1, msg_to_bit_it_8_vnu_30_in_2, msg_to_bit_it_8_vnu_31_in_0, msg_to_bit_it_8_vnu_31_in_1, msg_to_bit_it_8_vnu_31_in_2, msg_to_bit_it_8_vnu_32_in_0, msg_to_bit_it_8_vnu_32_in_1, msg_to_bit_it_8_vnu_32_in_2, msg_to_bit_it_8_vnu_33_in_0, msg_to_bit_it_8_vnu_33_in_1, msg_to_bit_it_8_vnu_33_in_2, msg_to_bit_it_8_vnu_34_in_0, msg_to_bit_it_8_vnu_34_in_1, msg_to_bit_it_8_vnu_34_in_2, msg_to_bit_it_8_vnu_35_in_0, msg_to_bit_it_8_vnu_35_in_1, msg_to_bit_it_8_vnu_35_in_2, msg_to_bit_it_8_vnu_36_in_0, msg_to_bit_it_8_vnu_36_in_1, msg_to_bit_it_8_vnu_36_in_2, msg_to_bit_it_8_vnu_37_in_0, msg_to_bit_it_8_vnu_37_in_1, msg_to_bit_it_8_vnu_37_in_2, msg_to_bit_it_8_vnu_38_in_0, msg_to_bit_it_8_vnu_38_in_1, msg_to_bit_it_8_vnu_38_in_2, msg_to_bit_it_8_vnu_39_in_0, msg_to_bit_it_8_vnu_39_in_1, msg_to_bit_it_8_vnu_39_in_2, msg_to_bit_it_8_vnu_40_in_0, msg_to_bit_it_8_vnu_40_in_1, msg_to_bit_it_8_vnu_40_in_2, msg_to_bit_it_8_vnu_41_in_0, msg_to_bit_it_8_vnu_41_in_1, msg_to_bit_it_8_vnu_41_in_2, msg_to_bit_it_8_vnu_42_in_0, msg_to_bit_it_8_vnu_42_in_1, msg_to_bit_it_8_vnu_42_in_2, msg_to_bit_it_8_vnu_43_in_0, msg_to_bit_it_8_vnu_43_in_1, msg_to_bit_it_8_vnu_43_in_2, msg_to_bit_it_8_vnu_44_in_0, msg_to_bit_it_8_vnu_44_in_1, msg_to_bit_it_8_vnu_44_in_2, msg_to_bit_it_8_vnu_45_in_0, msg_to_bit_it_8_vnu_45_in_1, msg_to_bit_it_8_vnu_45_in_2, msg_to_bit_it_8_vnu_46_in_0, msg_to_bit_it_8_vnu_46_in_1, msg_to_bit_it_8_vnu_46_in_2, msg_to_bit_it_8_vnu_47_in_0, msg_to_bit_it_8_vnu_47_in_1, msg_to_bit_it_8_vnu_47_in_2, msg_to_bit_it_8_vnu_48_in_0, msg_to_bit_it_8_vnu_48_in_1, msg_to_bit_it_8_vnu_48_in_2, msg_to_bit_it_8_vnu_49_in_0, msg_to_bit_it_8_vnu_49_in_1, msg_to_bit_it_8_vnu_49_in_2, msg_to_bit_it_8_vnu_50_in_0, msg_to_bit_it_8_vnu_50_in_1, msg_to_bit_it_8_vnu_50_in_2, msg_to_bit_it_8_vnu_51_in_0, msg_to_bit_it_8_vnu_51_in_1, msg_to_bit_it_8_vnu_51_in_2, msg_to_bit_it_8_vnu_52_in_0, msg_to_bit_it_8_vnu_52_in_1, msg_to_bit_it_8_vnu_52_in_2, msg_to_bit_it_8_vnu_53_in_0, msg_to_bit_it_8_vnu_53_in_1, msg_to_bit_it_8_vnu_53_in_2, msg_to_bit_it_8_vnu_54_in_0, msg_to_bit_it_8_vnu_54_in_1, msg_to_bit_it_8_vnu_54_in_2, msg_to_bit_it_8_vnu_55_in_0, msg_to_bit_it_8_vnu_55_in_1, msg_to_bit_it_8_vnu_55_in_2, msg_to_bit_it_8_vnu_56_in_0, msg_to_bit_it_8_vnu_56_in_1, msg_to_bit_it_8_vnu_56_in_2, msg_to_bit_it_8_vnu_57_in_0, msg_to_bit_it_8_vnu_57_in_1, msg_to_bit_it_8_vnu_57_in_2, msg_to_bit_it_8_vnu_58_in_0, msg_to_bit_it_8_vnu_58_in_1, msg_to_bit_it_8_vnu_58_in_2, msg_to_bit_it_8_vnu_59_in_0, msg_to_bit_it_8_vnu_59_in_1, msg_to_bit_it_8_vnu_59_in_2, msg_to_bit_it_8_vnu_60_in_0, msg_to_bit_it_8_vnu_60_in_1, msg_to_bit_it_8_vnu_60_in_2, msg_to_bit_it_8_vnu_61_in_0, msg_to_bit_it_8_vnu_61_in_1, msg_to_bit_it_8_vnu_61_in_2, msg_to_bit_it_8_vnu_62_in_0, msg_to_bit_it_8_vnu_62_in_1, msg_to_bit_it_8_vnu_62_in_2, msg_to_bit_it_8_vnu_63_in_0, msg_to_bit_it_8_vnu_63_in_1, msg_to_bit_it_8_vnu_63_in_2, msg_to_bit_it_8_vnu_64_in_0, msg_to_bit_it_8_vnu_64_in_1, msg_to_bit_it_8_vnu_64_in_2, msg_to_bit_it_8_vnu_65_in_0, msg_to_bit_it_8_vnu_65_in_1, msg_to_bit_it_8_vnu_65_in_2, msg_to_bit_it_8_vnu_66_in_0, msg_to_bit_it_8_vnu_66_in_1, msg_to_bit_it_8_vnu_66_in_2, msg_to_bit_it_8_vnu_67_in_0, msg_to_bit_it_8_vnu_67_in_1, msg_to_bit_it_8_vnu_67_in_2, msg_to_bit_it_8_vnu_68_in_0, msg_to_bit_it_8_vnu_68_in_1, msg_to_bit_it_8_vnu_68_in_2, msg_to_bit_it_8_vnu_69_in_0, msg_to_bit_it_8_vnu_69_in_1, msg_to_bit_it_8_vnu_69_in_2, msg_to_bit_it_8_vnu_70_in_0, msg_to_bit_it_8_vnu_70_in_1, msg_to_bit_it_8_vnu_70_in_2, msg_to_bit_it_8_vnu_71_in_0, msg_to_bit_it_8_vnu_71_in_1, msg_to_bit_it_8_vnu_71_in_2, msg_to_bit_it_8_vnu_72_in_0, msg_to_bit_it_8_vnu_72_in_1, msg_to_bit_it_8_vnu_72_in_2, msg_to_bit_it_8_vnu_73_in_0, msg_to_bit_it_8_vnu_73_in_1, msg_to_bit_it_8_vnu_73_in_2, msg_to_bit_it_8_vnu_74_in_0, msg_to_bit_it_8_vnu_74_in_1, msg_to_bit_it_8_vnu_74_in_2, msg_to_bit_it_8_vnu_75_in_0, msg_to_bit_it_8_vnu_75_in_1, msg_to_bit_it_8_vnu_75_in_2, msg_to_bit_it_8_vnu_76_in_0, msg_to_bit_it_8_vnu_76_in_1, msg_to_bit_it_8_vnu_76_in_2, msg_to_bit_it_8_vnu_77_in_0, msg_to_bit_it_8_vnu_77_in_1, msg_to_bit_it_8_vnu_77_in_2, msg_to_bit_it_8_vnu_78_in_0, msg_to_bit_it_8_vnu_78_in_1, msg_to_bit_it_8_vnu_78_in_2, msg_to_bit_it_8_vnu_79_in_0, msg_to_bit_it_8_vnu_79_in_1, msg_to_bit_it_8_vnu_79_in_2, msg_to_bit_it_8_vnu_80_in_0, msg_to_bit_it_8_vnu_80_in_1, msg_to_bit_it_8_vnu_80_in_2, msg_to_bit_it_8_vnu_81_in_0, msg_to_bit_it_8_vnu_81_in_1, msg_to_bit_it_8_vnu_81_in_2, msg_to_bit_it_8_vnu_82_in_0, msg_to_bit_it_8_vnu_82_in_1, msg_to_bit_it_8_vnu_82_in_2, msg_to_bit_it_8_vnu_83_in_0, msg_to_bit_it_8_vnu_83_in_1, msg_to_bit_it_8_vnu_83_in_2, msg_to_bit_it_8_vnu_84_in_0, msg_to_bit_it_8_vnu_84_in_1, msg_to_bit_it_8_vnu_84_in_2, msg_to_bit_it_8_vnu_85_in_0, msg_to_bit_it_8_vnu_85_in_1, msg_to_bit_it_8_vnu_85_in_2, msg_to_bit_it_8_vnu_86_in_0, msg_to_bit_it_8_vnu_86_in_1, msg_to_bit_it_8_vnu_86_in_2, msg_to_bit_it_8_vnu_87_in_0, msg_to_bit_it_8_vnu_87_in_1, msg_to_bit_it_8_vnu_87_in_2, msg_to_bit_it_8_vnu_88_in_0, msg_to_bit_it_8_vnu_88_in_1, msg_to_bit_it_8_vnu_88_in_2, msg_to_bit_it_8_vnu_89_in_0, msg_to_bit_it_8_vnu_89_in_1, msg_to_bit_it_8_vnu_89_in_2, msg_to_bit_it_8_vnu_90_in_0, msg_to_bit_it_8_vnu_90_in_1, msg_to_bit_it_8_vnu_90_in_2, msg_to_bit_it_8_vnu_91_in_0, msg_to_bit_it_8_vnu_91_in_1, msg_to_bit_it_8_vnu_91_in_2, msg_to_bit_it_8_vnu_92_in_0, msg_to_bit_it_8_vnu_92_in_1, msg_to_bit_it_8_vnu_92_in_2, msg_to_bit_it_8_vnu_93_in_0, msg_to_bit_it_8_vnu_93_in_1, msg_to_bit_it_8_vnu_93_in_2, msg_to_bit_it_8_vnu_94_in_0, msg_to_bit_it_8_vnu_94_in_1, msg_to_bit_it_8_vnu_94_in_2, msg_to_bit_it_8_vnu_95_in_0, msg_to_bit_it_8_vnu_95_in_1, msg_to_bit_it_8_vnu_95_in_2, msg_to_bit_it_8_vnu_96_in_0, msg_to_bit_it_8_vnu_96_in_1, msg_to_bit_it_8_vnu_96_in_2, msg_to_bit_it_8_vnu_97_in_0, msg_to_bit_it_8_vnu_97_in_1, msg_to_bit_it_8_vnu_97_in_2, msg_to_bit_it_8_vnu_98_in_0, msg_to_bit_it_8_vnu_98_in_1, msg_to_bit_it_8_vnu_98_in_2, msg_to_bit_it_8_vnu_99_in_0, msg_to_bit_it_8_vnu_99_in_1, msg_to_bit_it_8_vnu_99_in_2, msg_to_bit_it_8_vnu_100_in_0, msg_to_bit_it_8_vnu_100_in_1, msg_to_bit_it_8_vnu_100_in_2, msg_to_bit_it_8_vnu_101_in_0, msg_to_bit_it_8_vnu_101_in_1, msg_to_bit_it_8_vnu_101_in_2, msg_to_bit_it_8_vnu_102_in_0, msg_to_bit_it_8_vnu_102_in_1, msg_to_bit_it_8_vnu_102_in_2, msg_to_bit_it_8_vnu_103_in_0, msg_to_bit_it_8_vnu_103_in_1, msg_to_bit_it_8_vnu_103_in_2, msg_to_bit_it_8_vnu_104_in_0, msg_to_bit_it_8_vnu_104_in_1, msg_to_bit_it_8_vnu_104_in_2, msg_to_bit_it_8_vnu_105_in_0, msg_to_bit_it_8_vnu_105_in_1, msg_to_bit_it_8_vnu_105_in_2, msg_to_bit_it_8_vnu_106_in_0, msg_to_bit_it_8_vnu_106_in_1, msg_to_bit_it_8_vnu_106_in_2, msg_to_bit_it_8_vnu_107_in_0, msg_to_bit_it_8_vnu_107_in_1, msg_to_bit_it_8_vnu_107_in_2, msg_to_bit_it_8_vnu_108_in_0, msg_to_bit_it_8_vnu_108_in_1, msg_to_bit_it_8_vnu_108_in_2, msg_to_bit_it_8_vnu_109_in_0, msg_to_bit_it_8_vnu_109_in_1, msg_to_bit_it_8_vnu_109_in_2, msg_to_bit_it_8_vnu_110_in_0, msg_to_bit_it_8_vnu_110_in_1, msg_to_bit_it_8_vnu_110_in_2, msg_to_bit_it_8_vnu_111_in_0, msg_to_bit_it_8_vnu_111_in_1, msg_to_bit_it_8_vnu_111_in_2, msg_to_bit_it_8_vnu_112_in_0, msg_to_bit_it_8_vnu_112_in_1, msg_to_bit_it_8_vnu_112_in_2, msg_to_bit_it_8_vnu_113_in_0, msg_to_bit_it_8_vnu_113_in_1, msg_to_bit_it_8_vnu_113_in_2, msg_to_bit_it_8_vnu_114_in_0, msg_to_bit_it_8_vnu_114_in_1, msg_to_bit_it_8_vnu_114_in_2, msg_to_bit_it_8_vnu_115_in_0, msg_to_bit_it_8_vnu_115_in_1, msg_to_bit_it_8_vnu_115_in_2, msg_to_bit_it_8_vnu_116_in_0, msg_to_bit_it_8_vnu_116_in_1, msg_to_bit_it_8_vnu_116_in_2, msg_to_bit_it_8_vnu_117_in_0, msg_to_bit_it_8_vnu_117_in_1, msg_to_bit_it_8_vnu_117_in_2, msg_to_bit_it_8_vnu_118_in_0, msg_to_bit_it_8_vnu_118_in_1, msg_to_bit_it_8_vnu_118_in_2, msg_to_bit_it_8_vnu_119_in_0, msg_to_bit_it_8_vnu_119_in_1, msg_to_bit_it_8_vnu_119_in_2, msg_to_bit_it_8_vnu_120_in_0, msg_to_bit_it_8_vnu_120_in_1, msg_to_bit_it_8_vnu_120_in_2, msg_to_bit_it_8_vnu_121_in_0, msg_to_bit_it_8_vnu_121_in_1, msg_to_bit_it_8_vnu_121_in_2, msg_to_bit_it_8_vnu_122_in_0, msg_to_bit_it_8_vnu_122_in_1, msg_to_bit_it_8_vnu_122_in_2, msg_to_bit_it_8_vnu_123_in_0, msg_to_bit_it_8_vnu_123_in_1, msg_to_bit_it_8_vnu_123_in_2, msg_to_bit_it_8_vnu_124_in_0, msg_to_bit_it_8_vnu_124_in_1, msg_to_bit_it_8_vnu_124_in_2, msg_to_bit_it_8_vnu_125_in_0, msg_to_bit_it_8_vnu_125_in_1, msg_to_bit_it_8_vnu_125_in_2, msg_to_bit_it_8_vnu_126_in_0, msg_to_bit_it_8_vnu_126_in_1, msg_to_bit_it_8_vnu_126_in_2, msg_to_bit_it_8_vnu_127_in_0, msg_to_bit_it_8_vnu_127_in_1, msg_to_bit_it_8_vnu_127_in_2, msg_to_bit_it_8_vnu_128_in_0, msg_to_bit_it_8_vnu_128_in_1, msg_to_bit_it_8_vnu_128_in_2, msg_to_bit_it_8_vnu_129_in_0, msg_to_bit_it_8_vnu_129_in_1, msg_to_bit_it_8_vnu_129_in_2, msg_to_bit_it_8_vnu_130_in_0, msg_to_bit_it_8_vnu_130_in_1, msg_to_bit_it_8_vnu_130_in_2, msg_to_bit_it_8_vnu_131_in_0, msg_to_bit_it_8_vnu_131_in_1, msg_to_bit_it_8_vnu_131_in_2, msg_to_bit_it_8_vnu_132_in_0, msg_to_bit_it_8_vnu_132_in_1, msg_to_bit_it_8_vnu_132_in_2, msg_to_bit_it_8_vnu_133_in_0, msg_to_bit_it_8_vnu_133_in_1, msg_to_bit_it_8_vnu_133_in_2, msg_to_bit_it_8_vnu_134_in_0, msg_to_bit_it_8_vnu_134_in_1, msg_to_bit_it_8_vnu_134_in_2, msg_to_bit_it_8_vnu_135_in_0, msg_to_bit_it_8_vnu_135_in_1, msg_to_bit_it_8_vnu_135_in_2, msg_to_bit_it_8_vnu_136_in_0, msg_to_bit_it_8_vnu_136_in_1, msg_to_bit_it_8_vnu_136_in_2, msg_to_bit_it_8_vnu_137_in_0, msg_to_bit_it_8_vnu_137_in_1, msg_to_bit_it_8_vnu_137_in_2, msg_to_bit_it_8_vnu_138_in_0, msg_to_bit_it_8_vnu_138_in_1, msg_to_bit_it_8_vnu_138_in_2, msg_to_bit_it_8_vnu_139_in_0, msg_to_bit_it_8_vnu_139_in_1, msg_to_bit_it_8_vnu_139_in_2, msg_to_bit_it_8_vnu_140_in_0, msg_to_bit_it_8_vnu_140_in_1, msg_to_bit_it_8_vnu_140_in_2, msg_to_bit_it_8_vnu_141_in_0, msg_to_bit_it_8_vnu_141_in_1, msg_to_bit_it_8_vnu_141_in_2, msg_to_bit_it_8_vnu_142_in_0, msg_to_bit_it_8_vnu_142_in_1, msg_to_bit_it_8_vnu_142_in_2, msg_to_bit_it_8_vnu_143_in_0, msg_to_bit_it_8_vnu_143_in_1, msg_to_bit_it_8_vnu_143_in_2, msg_to_bit_it_8_vnu_144_in_0, msg_to_bit_it_8_vnu_144_in_1, msg_to_bit_it_8_vnu_144_in_2, msg_to_bit_it_8_vnu_145_in_0, msg_to_bit_it_8_vnu_145_in_1, msg_to_bit_it_8_vnu_145_in_2, msg_to_bit_it_8_vnu_146_in_0, msg_to_bit_it_8_vnu_146_in_1, msg_to_bit_it_8_vnu_146_in_2, msg_to_bit_it_8_vnu_147_in_0, msg_to_bit_it_8_vnu_147_in_1, msg_to_bit_it_8_vnu_147_in_2, msg_to_bit_it_8_vnu_148_in_0, msg_to_bit_it_8_vnu_148_in_1, msg_to_bit_it_8_vnu_148_in_2, msg_to_bit_it_8_vnu_149_in_0, msg_to_bit_it_8_vnu_149_in_1, msg_to_bit_it_8_vnu_149_in_2, msg_to_bit_it_8_vnu_150_in_0, msg_to_bit_it_8_vnu_150_in_1, msg_to_bit_it_8_vnu_150_in_2, msg_to_bit_it_8_vnu_151_in_0, msg_to_bit_it_8_vnu_151_in_1, msg_to_bit_it_8_vnu_151_in_2, msg_to_bit_it_8_vnu_152_in_0, msg_to_bit_it_8_vnu_152_in_1, msg_to_bit_it_8_vnu_152_in_2, msg_to_bit_it_8_vnu_153_in_0, msg_to_bit_it_8_vnu_153_in_1, msg_to_bit_it_8_vnu_153_in_2, msg_to_bit_it_8_vnu_154_in_0, msg_to_bit_it_8_vnu_154_in_1, msg_to_bit_it_8_vnu_154_in_2, msg_to_bit_it_8_vnu_155_in_0, msg_to_bit_it_8_vnu_155_in_1, msg_to_bit_it_8_vnu_155_in_2, msg_to_bit_it_8_vnu_156_in_0, msg_to_bit_it_8_vnu_156_in_1, msg_to_bit_it_8_vnu_156_in_2, msg_to_bit_it_8_vnu_157_in_0, msg_to_bit_it_8_vnu_157_in_1, msg_to_bit_it_8_vnu_157_in_2, msg_to_bit_it_8_vnu_158_in_0, msg_to_bit_it_8_vnu_158_in_1, msg_to_bit_it_8_vnu_158_in_2, msg_to_bit_it_8_vnu_159_in_0, msg_to_bit_it_8_vnu_159_in_1, msg_to_bit_it_8_vnu_159_in_2, msg_to_bit_it_8_vnu_160_in_0, msg_to_bit_it_8_vnu_160_in_1, msg_to_bit_it_8_vnu_160_in_2, msg_to_bit_it_8_vnu_161_in_0, msg_to_bit_it_8_vnu_161_in_1, msg_to_bit_it_8_vnu_161_in_2, msg_to_bit_it_8_vnu_162_in_0, msg_to_bit_it_8_vnu_162_in_1, msg_to_bit_it_8_vnu_162_in_2, msg_to_bit_it_8_vnu_163_in_0, msg_to_bit_it_8_vnu_163_in_1, msg_to_bit_it_8_vnu_163_in_2, msg_to_bit_it_8_vnu_164_in_0, msg_to_bit_it_8_vnu_164_in_1, msg_to_bit_it_8_vnu_164_in_2, msg_to_bit_it_8_vnu_165_in_0, msg_to_bit_it_8_vnu_165_in_1, msg_to_bit_it_8_vnu_165_in_2, msg_to_bit_it_8_vnu_166_in_0, msg_to_bit_it_8_vnu_166_in_1, msg_to_bit_it_8_vnu_166_in_2, msg_to_bit_it_8_vnu_167_in_0, msg_to_bit_it_8_vnu_167_in_1, msg_to_bit_it_8_vnu_167_in_2, msg_to_bit_it_8_vnu_168_in_0, msg_to_bit_it_8_vnu_168_in_1, msg_to_bit_it_8_vnu_168_in_2, msg_to_bit_it_8_vnu_169_in_0, msg_to_bit_it_8_vnu_169_in_1, msg_to_bit_it_8_vnu_169_in_2, msg_to_bit_it_8_vnu_170_in_0, msg_to_bit_it_8_vnu_170_in_1, msg_to_bit_it_8_vnu_170_in_2, msg_to_bit_it_8_vnu_171_in_0, msg_to_bit_it_8_vnu_171_in_1, msg_to_bit_it_8_vnu_171_in_2, msg_to_bit_it_8_vnu_172_in_0, msg_to_bit_it_8_vnu_172_in_1, msg_to_bit_it_8_vnu_172_in_2, msg_to_bit_it_8_vnu_173_in_0, msg_to_bit_it_8_vnu_173_in_1, msg_to_bit_it_8_vnu_173_in_2, msg_to_bit_it_8_vnu_174_in_0, msg_to_bit_it_8_vnu_174_in_1, msg_to_bit_it_8_vnu_174_in_2, msg_to_bit_it_8_vnu_175_in_0, msg_to_bit_it_8_vnu_175_in_1, msg_to_bit_it_8_vnu_175_in_2, msg_to_bit_it_8_vnu_176_in_0, msg_to_bit_it_8_vnu_176_in_1, msg_to_bit_it_8_vnu_176_in_2, msg_to_bit_it_8_vnu_177_in_0, msg_to_bit_it_8_vnu_177_in_1, msg_to_bit_it_8_vnu_177_in_2, msg_to_bit_it_8_vnu_178_in_0, msg_to_bit_it_8_vnu_178_in_1, msg_to_bit_it_8_vnu_178_in_2, msg_to_bit_it_8_vnu_179_in_0, msg_to_bit_it_8_vnu_179_in_1, msg_to_bit_it_8_vnu_179_in_2, msg_to_bit_it_8_vnu_180_in_0, msg_to_bit_it_8_vnu_180_in_1, msg_to_bit_it_8_vnu_180_in_2, msg_to_bit_it_8_vnu_181_in_0, msg_to_bit_it_8_vnu_181_in_1, msg_to_bit_it_8_vnu_181_in_2, msg_to_bit_it_8_vnu_182_in_0, msg_to_bit_it_8_vnu_182_in_1, msg_to_bit_it_8_vnu_182_in_2, msg_to_bit_it_8_vnu_183_in_0, msg_to_bit_it_8_vnu_183_in_1, msg_to_bit_it_8_vnu_183_in_2, msg_to_bit_it_8_vnu_184_in_0, msg_to_bit_it_8_vnu_184_in_1, msg_to_bit_it_8_vnu_184_in_2, msg_to_bit_it_8_vnu_185_in_0, msg_to_bit_it_8_vnu_185_in_1, msg_to_bit_it_8_vnu_185_in_2, msg_to_bit_it_8_vnu_186_in_0, msg_to_bit_it_8_vnu_186_in_1, msg_to_bit_it_8_vnu_186_in_2, msg_to_bit_it_8_vnu_187_in_0, msg_to_bit_it_8_vnu_187_in_1, msg_to_bit_it_8_vnu_187_in_2, msg_to_bit_it_8_vnu_188_in_0, msg_to_bit_it_8_vnu_188_in_1, msg_to_bit_it_8_vnu_188_in_2, msg_to_bit_it_8_vnu_189_in_0, msg_to_bit_it_8_vnu_189_in_1, msg_to_bit_it_8_vnu_189_in_2, msg_to_bit_it_8_vnu_190_in_0, msg_to_bit_it_8_vnu_190_in_1, msg_to_bit_it_8_vnu_190_in_2, msg_to_bit_it_8_vnu_191_in_0, msg_to_bit_it_8_vnu_191_in_1, msg_to_bit_it_8_vnu_191_in_2, msg_to_bit_it_8_vnu_192_in_0, msg_to_bit_it_8_vnu_192_in_1, msg_to_bit_it_8_vnu_192_in_2, msg_to_bit_it_8_vnu_193_in_0, msg_to_bit_it_8_vnu_193_in_1, msg_to_bit_it_8_vnu_193_in_2, msg_to_bit_it_8_vnu_194_in_0, msg_to_bit_it_8_vnu_194_in_1, msg_to_bit_it_8_vnu_194_in_2, msg_to_bit_it_8_vnu_195_in_0, msg_to_bit_it_8_vnu_195_in_1, msg_to_bit_it_8_vnu_195_in_2, msg_to_bit_it_8_vnu_196_in_0, msg_to_bit_it_8_vnu_196_in_1, msg_to_bit_it_8_vnu_196_in_2, msg_to_bit_it_8_vnu_197_in_0, msg_to_bit_it_8_vnu_197_in_1, msg_to_bit_it_8_vnu_197_in_2, msg_to_bit_it_9_vnu_0_in_0, msg_to_bit_it_9_vnu_0_in_1, msg_to_bit_it_9_vnu_0_in_2, msg_to_bit_it_9_vnu_1_in_0, msg_to_bit_it_9_vnu_1_in_1, msg_to_bit_it_9_vnu_1_in_2, msg_to_bit_it_9_vnu_2_in_0, msg_to_bit_it_9_vnu_2_in_1, msg_to_bit_it_9_vnu_2_in_2, msg_to_bit_it_9_vnu_3_in_0, msg_to_bit_it_9_vnu_3_in_1, msg_to_bit_it_9_vnu_3_in_2, msg_to_bit_it_9_vnu_4_in_0, msg_to_bit_it_9_vnu_4_in_1, msg_to_bit_it_9_vnu_4_in_2, msg_to_bit_it_9_vnu_5_in_0, msg_to_bit_it_9_vnu_5_in_1, msg_to_bit_it_9_vnu_5_in_2, msg_to_bit_it_9_vnu_6_in_0, msg_to_bit_it_9_vnu_6_in_1, msg_to_bit_it_9_vnu_6_in_2, msg_to_bit_it_9_vnu_7_in_0, msg_to_bit_it_9_vnu_7_in_1, msg_to_bit_it_9_vnu_7_in_2, msg_to_bit_it_9_vnu_8_in_0, msg_to_bit_it_9_vnu_8_in_1, msg_to_bit_it_9_vnu_8_in_2, msg_to_bit_it_9_vnu_9_in_0, msg_to_bit_it_9_vnu_9_in_1, msg_to_bit_it_9_vnu_9_in_2, msg_to_bit_it_9_vnu_10_in_0, msg_to_bit_it_9_vnu_10_in_1, msg_to_bit_it_9_vnu_10_in_2, msg_to_bit_it_9_vnu_11_in_0, msg_to_bit_it_9_vnu_11_in_1, msg_to_bit_it_9_vnu_11_in_2, msg_to_bit_it_9_vnu_12_in_0, msg_to_bit_it_9_vnu_12_in_1, msg_to_bit_it_9_vnu_12_in_2, msg_to_bit_it_9_vnu_13_in_0, msg_to_bit_it_9_vnu_13_in_1, msg_to_bit_it_9_vnu_13_in_2, msg_to_bit_it_9_vnu_14_in_0, msg_to_bit_it_9_vnu_14_in_1, msg_to_bit_it_9_vnu_14_in_2, msg_to_bit_it_9_vnu_15_in_0, msg_to_bit_it_9_vnu_15_in_1, msg_to_bit_it_9_vnu_15_in_2, msg_to_bit_it_9_vnu_16_in_0, msg_to_bit_it_9_vnu_16_in_1, msg_to_bit_it_9_vnu_16_in_2, msg_to_bit_it_9_vnu_17_in_0, msg_to_bit_it_9_vnu_17_in_1, msg_to_bit_it_9_vnu_17_in_2, msg_to_bit_it_9_vnu_18_in_0, msg_to_bit_it_9_vnu_18_in_1, msg_to_bit_it_9_vnu_18_in_2, msg_to_bit_it_9_vnu_19_in_0, msg_to_bit_it_9_vnu_19_in_1, msg_to_bit_it_9_vnu_19_in_2, msg_to_bit_it_9_vnu_20_in_0, msg_to_bit_it_9_vnu_20_in_1, msg_to_bit_it_9_vnu_20_in_2, msg_to_bit_it_9_vnu_21_in_0, msg_to_bit_it_9_vnu_21_in_1, msg_to_bit_it_9_vnu_21_in_2, msg_to_bit_it_9_vnu_22_in_0, msg_to_bit_it_9_vnu_22_in_1, msg_to_bit_it_9_vnu_22_in_2, msg_to_bit_it_9_vnu_23_in_0, msg_to_bit_it_9_vnu_23_in_1, msg_to_bit_it_9_vnu_23_in_2, msg_to_bit_it_9_vnu_24_in_0, msg_to_bit_it_9_vnu_24_in_1, msg_to_bit_it_9_vnu_24_in_2, msg_to_bit_it_9_vnu_25_in_0, msg_to_bit_it_9_vnu_25_in_1, msg_to_bit_it_9_vnu_25_in_2, msg_to_bit_it_9_vnu_26_in_0, msg_to_bit_it_9_vnu_26_in_1, msg_to_bit_it_9_vnu_26_in_2, msg_to_bit_it_9_vnu_27_in_0, msg_to_bit_it_9_vnu_27_in_1, msg_to_bit_it_9_vnu_27_in_2, msg_to_bit_it_9_vnu_28_in_0, msg_to_bit_it_9_vnu_28_in_1, msg_to_bit_it_9_vnu_28_in_2, msg_to_bit_it_9_vnu_29_in_0, msg_to_bit_it_9_vnu_29_in_1, msg_to_bit_it_9_vnu_29_in_2, msg_to_bit_it_9_vnu_30_in_0, msg_to_bit_it_9_vnu_30_in_1, msg_to_bit_it_9_vnu_30_in_2, msg_to_bit_it_9_vnu_31_in_0, msg_to_bit_it_9_vnu_31_in_1, msg_to_bit_it_9_vnu_31_in_2, msg_to_bit_it_9_vnu_32_in_0, msg_to_bit_it_9_vnu_32_in_1, msg_to_bit_it_9_vnu_32_in_2, msg_to_bit_it_9_vnu_33_in_0, msg_to_bit_it_9_vnu_33_in_1, msg_to_bit_it_9_vnu_33_in_2, msg_to_bit_it_9_vnu_34_in_0, msg_to_bit_it_9_vnu_34_in_1, msg_to_bit_it_9_vnu_34_in_2, msg_to_bit_it_9_vnu_35_in_0, msg_to_bit_it_9_vnu_35_in_1, msg_to_bit_it_9_vnu_35_in_2, msg_to_bit_it_9_vnu_36_in_0, msg_to_bit_it_9_vnu_36_in_1, msg_to_bit_it_9_vnu_36_in_2, msg_to_bit_it_9_vnu_37_in_0, msg_to_bit_it_9_vnu_37_in_1, msg_to_bit_it_9_vnu_37_in_2, msg_to_bit_it_9_vnu_38_in_0, msg_to_bit_it_9_vnu_38_in_1, msg_to_bit_it_9_vnu_38_in_2, msg_to_bit_it_9_vnu_39_in_0, msg_to_bit_it_9_vnu_39_in_1, msg_to_bit_it_9_vnu_39_in_2, msg_to_bit_it_9_vnu_40_in_0, msg_to_bit_it_9_vnu_40_in_1, msg_to_bit_it_9_vnu_40_in_2, msg_to_bit_it_9_vnu_41_in_0, msg_to_bit_it_9_vnu_41_in_1, msg_to_bit_it_9_vnu_41_in_2, msg_to_bit_it_9_vnu_42_in_0, msg_to_bit_it_9_vnu_42_in_1, msg_to_bit_it_9_vnu_42_in_2, msg_to_bit_it_9_vnu_43_in_0, msg_to_bit_it_9_vnu_43_in_1, msg_to_bit_it_9_vnu_43_in_2, msg_to_bit_it_9_vnu_44_in_0, msg_to_bit_it_9_vnu_44_in_1, msg_to_bit_it_9_vnu_44_in_2, msg_to_bit_it_9_vnu_45_in_0, msg_to_bit_it_9_vnu_45_in_1, msg_to_bit_it_9_vnu_45_in_2, msg_to_bit_it_9_vnu_46_in_0, msg_to_bit_it_9_vnu_46_in_1, msg_to_bit_it_9_vnu_46_in_2, msg_to_bit_it_9_vnu_47_in_0, msg_to_bit_it_9_vnu_47_in_1, msg_to_bit_it_9_vnu_47_in_2, msg_to_bit_it_9_vnu_48_in_0, msg_to_bit_it_9_vnu_48_in_1, msg_to_bit_it_9_vnu_48_in_2, msg_to_bit_it_9_vnu_49_in_0, msg_to_bit_it_9_vnu_49_in_1, msg_to_bit_it_9_vnu_49_in_2, msg_to_bit_it_9_vnu_50_in_0, msg_to_bit_it_9_vnu_50_in_1, msg_to_bit_it_9_vnu_50_in_2, msg_to_bit_it_9_vnu_51_in_0, msg_to_bit_it_9_vnu_51_in_1, msg_to_bit_it_9_vnu_51_in_2, msg_to_bit_it_9_vnu_52_in_0, msg_to_bit_it_9_vnu_52_in_1, msg_to_bit_it_9_vnu_52_in_2, msg_to_bit_it_9_vnu_53_in_0, msg_to_bit_it_9_vnu_53_in_1, msg_to_bit_it_9_vnu_53_in_2, msg_to_bit_it_9_vnu_54_in_0, msg_to_bit_it_9_vnu_54_in_1, msg_to_bit_it_9_vnu_54_in_2, msg_to_bit_it_9_vnu_55_in_0, msg_to_bit_it_9_vnu_55_in_1, msg_to_bit_it_9_vnu_55_in_2, msg_to_bit_it_9_vnu_56_in_0, msg_to_bit_it_9_vnu_56_in_1, msg_to_bit_it_9_vnu_56_in_2, msg_to_bit_it_9_vnu_57_in_0, msg_to_bit_it_9_vnu_57_in_1, msg_to_bit_it_9_vnu_57_in_2, msg_to_bit_it_9_vnu_58_in_0, msg_to_bit_it_9_vnu_58_in_1, msg_to_bit_it_9_vnu_58_in_2, msg_to_bit_it_9_vnu_59_in_0, msg_to_bit_it_9_vnu_59_in_1, msg_to_bit_it_9_vnu_59_in_2, msg_to_bit_it_9_vnu_60_in_0, msg_to_bit_it_9_vnu_60_in_1, msg_to_bit_it_9_vnu_60_in_2, msg_to_bit_it_9_vnu_61_in_0, msg_to_bit_it_9_vnu_61_in_1, msg_to_bit_it_9_vnu_61_in_2, msg_to_bit_it_9_vnu_62_in_0, msg_to_bit_it_9_vnu_62_in_1, msg_to_bit_it_9_vnu_62_in_2, msg_to_bit_it_9_vnu_63_in_0, msg_to_bit_it_9_vnu_63_in_1, msg_to_bit_it_9_vnu_63_in_2, msg_to_bit_it_9_vnu_64_in_0, msg_to_bit_it_9_vnu_64_in_1, msg_to_bit_it_9_vnu_64_in_2, msg_to_bit_it_9_vnu_65_in_0, msg_to_bit_it_9_vnu_65_in_1, msg_to_bit_it_9_vnu_65_in_2, msg_to_bit_it_9_vnu_66_in_0, msg_to_bit_it_9_vnu_66_in_1, msg_to_bit_it_9_vnu_66_in_2, msg_to_bit_it_9_vnu_67_in_0, msg_to_bit_it_9_vnu_67_in_1, msg_to_bit_it_9_vnu_67_in_2, msg_to_bit_it_9_vnu_68_in_0, msg_to_bit_it_9_vnu_68_in_1, msg_to_bit_it_9_vnu_68_in_2, msg_to_bit_it_9_vnu_69_in_0, msg_to_bit_it_9_vnu_69_in_1, msg_to_bit_it_9_vnu_69_in_2, msg_to_bit_it_9_vnu_70_in_0, msg_to_bit_it_9_vnu_70_in_1, msg_to_bit_it_9_vnu_70_in_2, msg_to_bit_it_9_vnu_71_in_0, msg_to_bit_it_9_vnu_71_in_1, msg_to_bit_it_9_vnu_71_in_2, msg_to_bit_it_9_vnu_72_in_0, msg_to_bit_it_9_vnu_72_in_1, msg_to_bit_it_9_vnu_72_in_2, msg_to_bit_it_9_vnu_73_in_0, msg_to_bit_it_9_vnu_73_in_1, msg_to_bit_it_9_vnu_73_in_2, msg_to_bit_it_9_vnu_74_in_0, msg_to_bit_it_9_vnu_74_in_1, msg_to_bit_it_9_vnu_74_in_2, msg_to_bit_it_9_vnu_75_in_0, msg_to_bit_it_9_vnu_75_in_1, msg_to_bit_it_9_vnu_75_in_2, msg_to_bit_it_9_vnu_76_in_0, msg_to_bit_it_9_vnu_76_in_1, msg_to_bit_it_9_vnu_76_in_2, msg_to_bit_it_9_vnu_77_in_0, msg_to_bit_it_9_vnu_77_in_1, msg_to_bit_it_9_vnu_77_in_2, msg_to_bit_it_9_vnu_78_in_0, msg_to_bit_it_9_vnu_78_in_1, msg_to_bit_it_9_vnu_78_in_2, msg_to_bit_it_9_vnu_79_in_0, msg_to_bit_it_9_vnu_79_in_1, msg_to_bit_it_9_vnu_79_in_2, msg_to_bit_it_9_vnu_80_in_0, msg_to_bit_it_9_vnu_80_in_1, msg_to_bit_it_9_vnu_80_in_2, msg_to_bit_it_9_vnu_81_in_0, msg_to_bit_it_9_vnu_81_in_1, msg_to_bit_it_9_vnu_81_in_2, msg_to_bit_it_9_vnu_82_in_0, msg_to_bit_it_9_vnu_82_in_1, msg_to_bit_it_9_vnu_82_in_2, msg_to_bit_it_9_vnu_83_in_0, msg_to_bit_it_9_vnu_83_in_1, msg_to_bit_it_9_vnu_83_in_2, msg_to_bit_it_9_vnu_84_in_0, msg_to_bit_it_9_vnu_84_in_1, msg_to_bit_it_9_vnu_84_in_2, msg_to_bit_it_9_vnu_85_in_0, msg_to_bit_it_9_vnu_85_in_1, msg_to_bit_it_9_vnu_85_in_2, msg_to_bit_it_9_vnu_86_in_0, msg_to_bit_it_9_vnu_86_in_1, msg_to_bit_it_9_vnu_86_in_2, msg_to_bit_it_9_vnu_87_in_0, msg_to_bit_it_9_vnu_87_in_1, msg_to_bit_it_9_vnu_87_in_2, msg_to_bit_it_9_vnu_88_in_0, msg_to_bit_it_9_vnu_88_in_1, msg_to_bit_it_9_vnu_88_in_2, msg_to_bit_it_9_vnu_89_in_0, msg_to_bit_it_9_vnu_89_in_1, msg_to_bit_it_9_vnu_89_in_2, msg_to_bit_it_9_vnu_90_in_0, msg_to_bit_it_9_vnu_90_in_1, msg_to_bit_it_9_vnu_90_in_2, msg_to_bit_it_9_vnu_91_in_0, msg_to_bit_it_9_vnu_91_in_1, msg_to_bit_it_9_vnu_91_in_2, msg_to_bit_it_9_vnu_92_in_0, msg_to_bit_it_9_vnu_92_in_1, msg_to_bit_it_9_vnu_92_in_2, msg_to_bit_it_9_vnu_93_in_0, msg_to_bit_it_9_vnu_93_in_1, msg_to_bit_it_9_vnu_93_in_2, msg_to_bit_it_9_vnu_94_in_0, msg_to_bit_it_9_vnu_94_in_1, msg_to_bit_it_9_vnu_94_in_2, msg_to_bit_it_9_vnu_95_in_0, msg_to_bit_it_9_vnu_95_in_1, msg_to_bit_it_9_vnu_95_in_2, msg_to_bit_it_9_vnu_96_in_0, msg_to_bit_it_9_vnu_96_in_1, msg_to_bit_it_9_vnu_96_in_2, msg_to_bit_it_9_vnu_97_in_0, msg_to_bit_it_9_vnu_97_in_1, msg_to_bit_it_9_vnu_97_in_2, msg_to_bit_it_9_vnu_98_in_0, msg_to_bit_it_9_vnu_98_in_1, msg_to_bit_it_9_vnu_98_in_2, msg_to_bit_it_9_vnu_99_in_0, msg_to_bit_it_9_vnu_99_in_1, msg_to_bit_it_9_vnu_99_in_2, msg_to_bit_it_9_vnu_100_in_0, msg_to_bit_it_9_vnu_100_in_1, msg_to_bit_it_9_vnu_100_in_2, msg_to_bit_it_9_vnu_101_in_0, msg_to_bit_it_9_vnu_101_in_1, msg_to_bit_it_9_vnu_101_in_2, msg_to_bit_it_9_vnu_102_in_0, msg_to_bit_it_9_vnu_102_in_1, msg_to_bit_it_9_vnu_102_in_2, msg_to_bit_it_9_vnu_103_in_0, msg_to_bit_it_9_vnu_103_in_1, msg_to_bit_it_9_vnu_103_in_2, msg_to_bit_it_9_vnu_104_in_0, msg_to_bit_it_9_vnu_104_in_1, msg_to_bit_it_9_vnu_104_in_2, msg_to_bit_it_9_vnu_105_in_0, msg_to_bit_it_9_vnu_105_in_1, msg_to_bit_it_9_vnu_105_in_2, msg_to_bit_it_9_vnu_106_in_0, msg_to_bit_it_9_vnu_106_in_1, msg_to_bit_it_9_vnu_106_in_2, msg_to_bit_it_9_vnu_107_in_0, msg_to_bit_it_9_vnu_107_in_1, msg_to_bit_it_9_vnu_107_in_2, msg_to_bit_it_9_vnu_108_in_0, msg_to_bit_it_9_vnu_108_in_1, msg_to_bit_it_9_vnu_108_in_2, msg_to_bit_it_9_vnu_109_in_0, msg_to_bit_it_9_vnu_109_in_1, msg_to_bit_it_9_vnu_109_in_2, msg_to_bit_it_9_vnu_110_in_0, msg_to_bit_it_9_vnu_110_in_1, msg_to_bit_it_9_vnu_110_in_2, msg_to_bit_it_9_vnu_111_in_0, msg_to_bit_it_9_vnu_111_in_1, msg_to_bit_it_9_vnu_111_in_2, msg_to_bit_it_9_vnu_112_in_0, msg_to_bit_it_9_vnu_112_in_1, msg_to_bit_it_9_vnu_112_in_2, msg_to_bit_it_9_vnu_113_in_0, msg_to_bit_it_9_vnu_113_in_1, msg_to_bit_it_9_vnu_113_in_2, msg_to_bit_it_9_vnu_114_in_0, msg_to_bit_it_9_vnu_114_in_1, msg_to_bit_it_9_vnu_114_in_2, msg_to_bit_it_9_vnu_115_in_0, msg_to_bit_it_9_vnu_115_in_1, msg_to_bit_it_9_vnu_115_in_2, msg_to_bit_it_9_vnu_116_in_0, msg_to_bit_it_9_vnu_116_in_1, msg_to_bit_it_9_vnu_116_in_2, msg_to_bit_it_9_vnu_117_in_0, msg_to_bit_it_9_vnu_117_in_1, msg_to_bit_it_9_vnu_117_in_2, msg_to_bit_it_9_vnu_118_in_0, msg_to_bit_it_9_vnu_118_in_1, msg_to_bit_it_9_vnu_118_in_2, msg_to_bit_it_9_vnu_119_in_0, msg_to_bit_it_9_vnu_119_in_1, msg_to_bit_it_9_vnu_119_in_2, msg_to_bit_it_9_vnu_120_in_0, msg_to_bit_it_9_vnu_120_in_1, msg_to_bit_it_9_vnu_120_in_2, msg_to_bit_it_9_vnu_121_in_0, msg_to_bit_it_9_vnu_121_in_1, msg_to_bit_it_9_vnu_121_in_2, msg_to_bit_it_9_vnu_122_in_0, msg_to_bit_it_9_vnu_122_in_1, msg_to_bit_it_9_vnu_122_in_2, msg_to_bit_it_9_vnu_123_in_0, msg_to_bit_it_9_vnu_123_in_1, msg_to_bit_it_9_vnu_123_in_2, msg_to_bit_it_9_vnu_124_in_0, msg_to_bit_it_9_vnu_124_in_1, msg_to_bit_it_9_vnu_124_in_2, msg_to_bit_it_9_vnu_125_in_0, msg_to_bit_it_9_vnu_125_in_1, msg_to_bit_it_9_vnu_125_in_2, msg_to_bit_it_9_vnu_126_in_0, msg_to_bit_it_9_vnu_126_in_1, msg_to_bit_it_9_vnu_126_in_2, msg_to_bit_it_9_vnu_127_in_0, msg_to_bit_it_9_vnu_127_in_1, msg_to_bit_it_9_vnu_127_in_2, msg_to_bit_it_9_vnu_128_in_0, msg_to_bit_it_9_vnu_128_in_1, msg_to_bit_it_9_vnu_128_in_2, msg_to_bit_it_9_vnu_129_in_0, msg_to_bit_it_9_vnu_129_in_1, msg_to_bit_it_9_vnu_129_in_2, msg_to_bit_it_9_vnu_130_in_0, msg_to_bit_it_9_vnu_130_in_1, msg_to_bit_it_9_vnu_130_in_2, msg_to_bit_it_9_vnu_131_in_0, msg_to_bit_it_9_vnu_131_in_1, msg_to_bit_it_9_vnu_131_in_2, msg_to_bit_it_9_vnu_132_in_0, msg_to_bit_it_9_vnu_132_in_1, msg_to_bit_it_9_vnu_132_in_2, msg_to_bit_it_9_vnu_133_in_0, msg_to_bit_it_9_vnu_133_in_1, msg_to_bit_it_9_vnu_133_in_2, msg_to_bit_it_9_vnu_134_in_0, msg_to_bit_it_9_vnu_134_in_1, msg_to_bit_it_9_vnu_134_in_2, msg_to_bit_it_9_vnu_135_in_0, msg_to_bit_it_9_vnu_135_in_1, msg_to_bit_it_9_vnu_135_in_2, msg_to_bit_it_9_vnu_136_in_0, msg_to_bit_it_9_vnu_136_in_1, msg_to_bit_it_9_vnu_136_in_2, msg_to_bit_it_9_vnu_137_in_0, msg_to_bit_it_9_vnu_137_in_1, msg_to_bit_it_9_vnu_137_in_2, msg_to_bit_it_9_vnu_138_in_0, msg_to_bit_it_9_vnu_138_in_1, msg_to_bit_it_9_vnu_138_in_2, msg_to_bit_it_9_vnu_139_in_0, msg_to_bit_it_9_vnu_139_in_1, msg_to_bit_it_9_vnu_139_in_2, msg_to_bit_it_9_vnu_140_in_0, msg_to_bit_it_9_vnu_140_in_1, msg_to_bit_it_9_vnu_140_in_2, msg_to_bit_it_9_vnu_141_in_0, msg_to_bit_it_9_vnu_141_in_1, msg_to_bit_it_9_vnu_141_in_2, msg_to_bit_it_9_vnu_142_in_0, msg_to_bit_it_9_vnu_142_in_1, msg_to_bit_it_9_vnu_142_in_2, msg_to_bit_it_9_vnu_143_in_0, msg_to_bit_it_9_vnu_143_in_1, msg_to_bit_it_9_vnu_143_in_2, msg_to_bit_it_9_vnu_144_in_0, msg_to_bit_it_9_vnu_144_in_1, msg_to_bit_it_9_vnu_144_in_2, msg_to_bit_it_9_vnu_145_in_0, msg_to_bit_it_9_vnu_145_in_1, msg_to_bit_it_9_vnu_145_in_2, msg_to_bit_it_9_vnu_146_in_0, msg_to_bit_it_9_vnu_146_in_1, msg_to_bit_it_9_vnu_146_in_2, msg_to_bit_it_9_vnu_147_in_0, msg_to_bit_it_9_vnu_147_in_1, msg_to_bit_it_9_vnu_147_in_2, msg_to_bit_it_9_vnu_148_in_0, msg_to_bit_it_9_vnu_148_in_1, msg_to_bit_it_9_vnu_148_in_2, msg_to_bit_it_9_vnu_149_in_0, msg_to_bit_it_9_vnu_149_in_1, msg_to_bit_it_9_vnu_149_in_2, msg_to_bit_it_9_vnu_150_in_0, msg_to_bit_it_9_vnu_150_in_1, msg_to_bit_it_9_vnu_150_in_2, msg_to_bit_it_9_vnu_151_in_0, msg_to_bit_it_9_vnu_151_in_1, msg_to_bit_it_9_vnu_151_in_2, msg_to_bit_it_9_vnu_152_in_0, msg_to_bit_it_9_vnu_152_in_1, msg_to_bit_it_9_vnu_152_in_2, msg_to_bit_it_9_vnu_153_in_0, msg_to_bit_it_9_vnu_153_in_1, msg_to_bit_it_9_vnu_153_in_2, msg_to_bit_it_9_vnu_154_in_0, msg_to_bit_it_9_vnu_154_in_1, msg_to_bit_it_9_vnu_154_in_2, msg_to_bit_it_9_vnu_155_in_0, msg_to_bit_it_9_vnu_155_in_1, msg_to_bit_it_9_vnu_155_in_2, msg_to_bit_it_9_vnu_156_in_0, msg_to_bit_it_9_vnu_156_in_1, msg_to_bit_it_9_vnu_156_in_2, msg_to_bit_it_9_vnu_157_in_0, msg_to_bit_it_9_vnu_157_in_1, msg_to_bit_it_9_vnu_157_in_2, msg_to_bit_it_9_vnu_158_in_0, msg_to_bit_it_9_vnu_158_in_1, msg_to_bit_it_9_vnu_158_in_2, msg_to_bit_it_9_vnu_159_in_0, msg_to_bit_it_9_vnu_159_in_1, msg_to_bit_it_9_vnu_159_in_2, msg_to_bit_it_9_vnu_160_in_0, msg_to_bit_it_9_vnu_160_in_1, msg_to_bit_it_9_vnu_160_in_2, msg_to_bit_it_9_vnu_161_in_0, msg_to_bit_it_9_vnu_161_in_1, msg_to_bit_it_9_vnu_161_in_2, msg_to_bit_it_9_vnu_162_in_0, msg_to_bit_it_9_vnu_162_in_1, msg_to_bit_it_9_vnu_162_in_2, msg_to_bit_it_9_vnu_163_in_0, msg_to_bit_it_9_vnu_163_in_1, msg_to_bit_it_9_vnu_163_in_2, msg_to_bit_it_9_vnu_164_in_0, msg_to_bit_it_9_vnu_164_in_1, msg_to_bit_it_9_vnu_164_in_2, msg_to_bit_it_9_vnu_165_in_0, msg_to_bit_it_9_vnu_165_in_1, msg_to_bit_it_9_vnu_165_in_2, msg_to_bit_it_9_vnu_166_in_0, msg_to_bit_it_9_vnu_166_in_1, msg_to_bit_it_9_vnu_166_in_2, msg_to_bit_it_9_vnu_167_in_0, msg_to_bit_it_9_vnu_167_in_1, msg_to_bit_it_9_vnu_167_in_2, msg_to_bit_it_9_vnu_168_in_0, msg_to_bit_it_9_vnu_168_in_1, msg_to_bit_it_9_vnu_168_in_2, msg_to_bit_it_9_vnu_169_in_0, msg_to_bit_it_9_vnu_169_in_1, msg_to_bit_it_9_vnu_169_in_2, msg_to_bit_it_9_vnu_170_in_0, msg_to_bit_it_9_vnu_170_in_1, msg_to_bit_it_9_vnu_170_in_2, msg_to_bit_it_9_vnu_171_in_0, msg_to_bit_it_9_vnu_171_in_1, msg_to_bit_it_9_vnu_171_in_2, msg_to_bit_it_9_vnu_172_in_0, msg_to_bit_it_9_vnu_172_in_1, msg_to_bit_it_9_vnu_172_in_2, msg_to_bit_it_9_vnu_173_in_0, msg_to_bit_it_9_vnu_173_in_1, msg_to_bit_it_9_vnu_173_in_2, msg_to_bit_it_9_vnu_174_in_0, msg_to_bit_it_9_vnu_174_in_1, msg_to_bit_it_9_vnu_174_in_2, msg_to_bit_it_9_vnu_175_in_0, msg_to_bit_it_9_vnu_175_in_1, msg_to_bit_it_9_vnu_175_in_2, msg_to_bit_it_9_vnu_176_in_0, msg_to_bit_it_9_vnu_176_in_1, msg_to_bit_it_9_vnu_176_in_2, msg_to_bit_it_9_vnu_177_in_0, msg_to_bit_it_9_vnu_177_in_1, msg_to_bit_it_9_vnu_177_in_2, msg_to_bit_it_9_vnu_178_in_0, msg_to_bit_it_9_vnu_178_in_1, msg_to_bit_it_9_vnu_178_in_2, msg_to_bit_it_9_vnu_179_in_0, msg_to_bit_it_9_vnu_179_in_1, msg_to_bit_it_9_vnu_179_in_2, msg_to_bit_it_9_vnu_180_in_0, msg_to_bit_it_9_vnu_180_in_1, msg_to_bit_it_9_vnu_180_in_2, msg_to_bit_it_9_vnu_181_in_0, msg_to_bit_it_9_vnu_181_in_1, msg_to_bit_it_9_vnu_181_in_2, msg_to_bit_it_9_vnu_182_in_0, msg_to_bit_it_9_vnu_182_in_1, msg_to_bit_it_9_vnu_182_in_2, msg_to_bit_it_9_vnu_183_in_0, msg_to_bit_it_9_vnu_183_in_1, msg_to_bit_it_9_vnu_183_in_2, msg_to_bit_it_9_vnu_184_in_0, msg_to_bit_it_9_vnu_184_in_1, msg_to_bit_it_9_vnu_184_in_2, msg_to_bit_it_9_vnu_185_in_0, msg_to_bit_it_9_vnu_185_in_1, msg_to_bit_it_9_vnu_185_in_2, msg_to_bit_it_9_vnu_186_in_0, msg_to_bit_it_9_vnu_186_in_1, msg_to_bit_it_9_vnu_186_in_2, msg_to_bit_it_9_vnu_187_in_0, msg_to_bit_it_9_vnu_187_in_1, msg_to_bit_it_9_vnu_187_in_2, msg_to_bit_it_9_vnu_188_in_0, msg_to_bit_it_9_vnu_188_in_1, msg_to_bit_it_9_vnu_188_in_2, msg_to_bit_it_9_vnu_189_in_0, msg_to_bit_it_9_vnu_189_in_1, msg_to_bit_it_9_vnu_189_in_2, msg_to_bit_it_9_vnu_190_in_0, msg_to_bit_it_9_vnu_190_in_1, msg_to_bit_it_9_vnu_190_in_2, msg_to_bit_it_9_vnu_191_in_0, msg_to_bit_it_9_vnu_191_in_1, msg_to_bit_it_9_vnu_191_in_2, msg_to_bit_it_9_vnu_192_in_0, msg_to_bit_it_9_vnu_192_in_1, msg_to_bit_it_9_vnu_192_in_2, msg_to_bit_it_9_vnu_193_in_0, msg_to_bit_it_9_vnu_193_in_1, msg_to_bit_it_9_vnu_193_in_2, msg_to_bit_it_9_vnu_194_in_0, msg_to_bit_it_9_vnu_194_in_1, msg_to_bit_it_9_vnu_194_in_2, msg_to_bit_it_9_vnu_195_in_0, msg_to_bit_it_9_vnu_195_in_1, msg_to_bit_it_9_vnu_195_in_2, msg_to_bit_it_9_vnu_196_in_0, msg_to_bit_it_9_vnu_196_in_1, msg_to_bit_it_9_vnu_196_in_2, msg_to_bit_it_9_vnu_197_in_0, msg_to_bit_it_9_vnu_197_in_1, msg_to_bit_it_9_vnu_197_in_2, msg_to_bit_it_10_vnu_0_in_0, msg_to_bit_it_10_vnu_0_in_1, msg_to_bit_it_10_vnu_0_in_2, msg_to_bit_it_10_vnu_1_in_0, msg_to_bit_it_10_vnu_1_in_1, msg_to_bit_it_10_vnu_1_in_2, msg_to_bit_it_10_vnu_2_in_0, msg_to_bit_it_10_vnu_2_in_1, msg_to_bit_it_10_vnu_2_in_2, msg_to_bit_it_10_vnu_3_in_0, msg_to_bit_it_10_vnu_3_in_1, msg_to_bit_it_10_vnu_3_in_2, msg_to_bit_it_10_vnu_4_in_0, msg_to_bit_it_10_vnu_4_in_1, msg_to_bit_it_10_vnu_4_in_2, msg_to_bit_it_10_vnu_5_in_0, msg_to_bit_it_10_vnu_5_in_1, msg_to_bit_it_10_vnu_5_in_2, msg_to_bit_it_10_vnu_6_in_0, msg_to_bit_it_10_vnu_6_in_1, msg_to_bit_it_10_vnu_6_in_2, msg_to_bit_it_10_vnu_7_in_0, msg_to_bit_it_10_vnu_7_in_1, msg_to_bit_it_10_vnu_7_in_2, msg_to_bit_it_10_vnu_8_in_0, msg_to_bit_it_10_vnu_8_in_1, msg_to_bit_it_10_vnu_8_in_2, msg_to_bit_it_10_vnu_9_in_0, msg_to_bit_it_10_vnu_9_in_1, msg_to_bit_it_10_vnu_9_in_2, msg_to_bit_it_10_vnu_10_in_0, msg_to_bit_it_10_vnu_10_in_1, msg_to_bit_it_10_vnu_10_in_2, msg_to_bit_it_10_vnu_11_in_0, msg_to_bit_it_10_vnu_11_in_1, msg_to_bit_it_10_vnu_11_in_2, msg_to_bit_it_10_vnu_12_in_0, msg_to_bit_it_10_vnu_12_in_1, msg_to_bit_it_10_vnu_12_in_2, msg_to_bit_it_10_vnu_13_in_0, msg_to_bit_it_10_vnu_13_in_1, msg_to_bit_it_10_vnu_13_in_2, msg_to_bit_it_10_vnu_14_in_0, msg_to_bit_it_10_vnu_14_in_1, msg_to_bit_it_10_vnu_14_in_2, msg_to_bit_it_10_vnu_15_in_0, msg_to_bit_it_10_vnu_15_in_1, msg_to_bit_it_10_vnu_15_in_2, msg_to_bit_it_10_vnu_16_in_0, msg_to_bit_it_10_vnu_16_in_1, msg_to_bit_it_10_vnu_16_in_2, msg_to_bit_it_10_vnu_17_in_0, msg_to_bit_it_10_vnu_17_in_1, msg_to_bit_it_10_vnu_17_in_2, msg_to_bit_it_10_vnu_18_in_0, msg_to_bit_it_10_vnu_18_in_1, msg_to_bit_it_10_vnu_18_in_2, msg_to_bit_it_10_vnu_19_in_0, msg_to_bit_it_10_vnu_19_in_1, msg_to_bit_it_10_vnu_19_in_2, msg_to_bit_it_10_vnu_20_in_0, msg_to_bit_it_10_vnu_20_in_1, msg_to_bit_it_10_vnu_20_in_2, msg_to_bit_it_10_vnu_21_in_0, msg_to_bit_it_10_vnu_21_in_1, msg_to_bit_it_10_vnu_21_in_2, msg_to_bit_it_10_vnu_22_in_0, msg_to_bit_it_10_vnu_22_in_1, msg_to_bit_it_10_vnu_22_in_2, msg_to_bit_it_10_vnu_23_in_0, msg_to_bit_it_10_vnu_23_in_1, msg_to_bit_it_10_vnu_23_in_2, msg_to_bit_it_10_vnu_24_in_0, msg_to_bit_it_10_vnu_24_in_1, msg_to_bit_it_10_vnu_24_in_2, msg_to_bit_it_10_vnu_25_in_0, msg_to_bit_it_10_vnu_25_in_1, msg_to_bit_it_10_vnu_25_in_2, msg_to_bit_it_10_vnu_26_in_0, msg_to_bit_it_10_vnu_26_in_1, msg_to_bit_it_10_vnu_26_in_2, msg_to_bit_it_10_vnu_27_in_0, msg_to_bit_it_10_vnu_27_in_1, msg_to_bit_it_10_vnu_27_in_2, msg_to_bit_it_10_vnu_28_in_0, msg_to_bit_it_10_vnu_28_in_1, msg_to_bit_it_10_vnu_28_in_2, msg_to_bit_it_10_vnu_29_in_0, msg_to_bit_it_10_vnu_29_in_1, msg_to_bit_it_10_vnu_29_in_2, msg_to_bit_it_10_vnu_30_in_0, msg_to_bit_it_10_vnu_30_in_1, msg_to_bit_it_10_vnu_30_in_2, msg_to_bit_it_10_vnu_31_in_0, msg_to_bit_it_10_vnu_31_in_1, msg_to_bit_it_10_vnu_31_in_2, msg_to_bit_it_10_vnu_32_in_0, msg_to_bit_it_10_vnu_32_in_1, msg_to_bit_it_10_vnu_32_in_2, msg_to_bit_it_10_vnu_33_in_0, msg_to_bit_it_10_vnu_33_in_1, msg_to_bit_it_10_vnu_33_in_2, msg_to_bit_it_10_vnu_34_in_0, msg_to_bit_it_10_vnu_34_in_1, msg_to_bit_it_10_vnu_34_in_2, msg_to_bit_it_10_vnu_35_in_0, msg_to_bit_it_10_vnu_35_in_1, msg_to_bit_it_10_vnu_35_in_2, msg_to_bit_it_10_vnu_36_in_0, msg_to_bit_it_10_vnu_36_in_1, msg_to_bit_it_10_vnu_36_in_2, msg_to_bit_it_10_vnu_37_in_0, msg_to_bit_it_10_vnu_37_in_1, msg_to_bit_it_10_vnu_37_in_2, msg_to_bit_it_10_vnu_38_in_0, msg_to_bit_it_10_vnu_38_in_1, msg_to_bit_it_10_vnu_38_in_2, msg_to_bit_it_10_vnu_39_in_0, msg_to_bit_it_10_vnu_39_in_1, msg_to_bit_it_10_vnu_39_in_2, msg_to_bit_it_10_vnu_40_in_0, msg_to_bit_it_10_vnu_40_in_1, msg_to_bit_it_10_vnu_40_in_2, msg_to_bit_it_10_vnu_41_in_0, msg_to_bit_it_10_vnu_41_in_1, msg_to_bit_it_10_vnu_41_in_2, msg_to_bit_it_10_vnu_42_in_0, msg_to_bit_it_10_vnu_42_in_1, msg_to_bit_it_10_vnu_42_in_2, msg_to_bit_it_10_vnu_43_in_0, msg_to_bit_it_10_vnu_43_in_1, msg_to_bit_it_10_vnu_43_in_2, msg_to_bit_it_10_vnu_44_in_0, msg_to_bit_it_10_vnu_44_in_1, msg_to_bit_it_10_vnu_44_in_2, msg_to_bit_it_10_vnu_45_in_0, msg_to_bit_it_10_vnu_45_in_1, msg_to_bit_it_10_vnu_45_in_2, msg_to_bit_it_10_vnu_46_in_0, msg_to_bit_it_10_vnu_46_in_1, msg_to_bit_it_10_vnu_46_in_2, msg_to_bit_it_10_vnu_47_in_0, msg_to_bit_it_10_vnu_47_in_1, msg_to_bit_it_10_vnu_47_in_2, msg_to_bit_it_10_vnu_48_in_0, msg_to_bit_it_10_vnu_48_in_1, msg_to_bit_it_10_vnu_48_in_2, msg_to_bit_it_10_vnu_49_in_0, msg_to_bit_it_10_vnu_49_in_1, msg_to_bit_it_10_vnu_49_in_2, msg_to_bit_it_10_vnu_50_in_0, msg_to_bit_it_10_vnu_50_in_1, msg_to_bit_it_10_vnu_50_in_2, msg_to_bit_it_10_vnu_51_in_0, msg_to_bit_it_10_vnu_51_in_1, msg_to_bit_it_10_vnu_51_in_2, msg_to_bit_it_10_vnu_52_in_0, msg_to_bit_it_10_vnu_52_in_1, msg_to_bit_it_10_vnu_52_in_2, msg_to_bit_it_10_vnu_53_in_0, msg_to_bit_it_10_vnu_53_in_1, msg_to_bit_it_10_vnu_53_in_2, msg_to_bit_it_10_vnu_54_in_0, msg_to_bit_it_10_vnu_54_in_1, msg_to_bit_it_10_vnu_54_in_2, msg_to_bit_it_10_vnu_55_in_0, msg_to_bit_it_10_vnu_55_in_1, msg_to_bit_it_10_vnu_55_in_2, msg_to_bit_it_10_vnu_56_in_0, msg_to_bit_it_10_vnu_56_in_1, msg_to_bit_it_10_vnu_56_in_2, msg_to_bit_it_10_vnu_57_in_0, msg_to_bit_it_10_vnu_57_in_1, msg_to_bit_it_10_vnu_57_in_2, msg_to_bit_it_10_vnu_58_in_0, msg_to_bit_it_10_vnu_58_in_1, msg_to_bit_it_10_vnu_58_in_2, msg_to_bit_it_10_vnu_59_in_0, msg_to_bit_it_10_vnu_59_in_1, msg_to_bit_it_10_vnu_59_in_2, msg_to_bit_it_10_vnu_60_in_0, msg_to_bit_it_10_vnu_60_in_1, msg_to_bit_it_10_vnu_60_in_2, msg_to_bit_it_10_vnu_61_in_0, msg_to_bit_it_10_vnu_61_in_1, msg_to_bit_it_10_vnu_61_in_2, msg_to_bit_it_10_vnu_62_in_0, msg_to_bit_it_10_vnu_62_in_1, msg_to_bit_it_10_vnu_62_in_2, msg_to_bit_it_10_vnu_63_in_0, msg_to_bit_it_10_vnu_63_in_1, msg_to_bit_it_10_vnu_63_in_2, msg_to_bit_it_10_vnu_64_in_0, msg_to_bit_it_10_vnu_64_in_1, msg_to_bit_it_10_vnu_64_in_2, msg_to_bit_it_10_vnu_65_in_0, msg_to_bit_it_10_vnu_65_in_1, msg_to_bit_it_10_vnu_65_in_2, msg_to_bit_it_10_vnu_66_in_0, msg_to_bit_it_10_vnu_66_in_1, msg_to_bit_it_10_vnu_66_in_2, msg_to_bit_it_10_vnu_67_in_0, msg_to_bit_it_10_vnu_67_in_1, msg_to_bit_it_10_vnu_67_in_2, msg_to_bit_it_10_vnu_68_in_0, msg_to_bit_it_10_vnu_68_in_1, msg_to_bit_it_10_vnu_68_in_2, msg_to_bit_it_10_vnu_69_in_0, msg_to_bit_it_10_vnu_69_in_1, msg_to_bit_it_10_vnu_69_in_2, msg_to_bit_it_10_vnu_70_in_0, msg_to_bit_it_10_vnu_70_in_1, msg_to_bit_it_10_vnu_70_in_2, msg_to_bit_it_10_vnu_71_in_0, msg_to_bit_it_10_vnu_71_in_1, msg_to_bit_it_10_vnu_71_in_2, msg_to_bit_it_10_vnu_72_in_0, msg_to_bit_it_10_vnu_72_in_1, msg_to_bit_it_10_vnu_72_in_2, msg_to_bit_it_10_vnu_73_in_0, msg_to_bit_it_10_vnu_73_in_1, msg_to_bit_it_10_vnu_73_in_2, msg_to_bit_it_10_vnu_74_in_0, msg_to_bit_it_10_vnu_74_in_1, msg_to_bit_it_10_vnu_74_in_2, msg_to_bit_it_10_vnu_75_in_0, msg_to_bit_it_10_vnu_75_in_1, msg_to_bit_it_10_vnu_75_in_2, msg_to_bit_it_10_vnu_76_in_0, msg_to_bit_it_10_vnu_76_in_1, msg_to_bit_it_10_vnu_76_in_2, msg_to_bit_it_10_vnu_77_in_0, msg_to_bit_it_10_vnu_77_in_1, msg_to_bit_it_10_vnu_77_in_2, msg_to_bit_it_10_vnu_78_in_0, msg_to_bit_it_10_vnu_78_in_1, msg_to_bit_it_10_vnu_78_in_2, msg_to_bit_it_10_vnu_79_in_0, msg_to_bit_it_10_vnu_79_in_1, msg_to_bit_it_10_vnu_79_in_2, msg_to_bit_it_10_vnu_80_in_0, msg_to_bit_it_10_vnu_80_in_1, msg_to_bit_it_10_vnu_80_in_2, msg_to_bit_it_10_vnu_81_in_0, msg_to_bit_it_10_vnu_81_in_1, msg_to_bit_it_10_vnu_81_in_2, msg_to_bit_it_10_vnu_82_in_0, msg_to_bit_it_10_vnu_82_in_1, msg_to_bit_it_10_vnu_82_in_2, msg_to_bit_it_10_vnu_83_in_0, msg_to_bit_it_10_vnu_83_in_1, msg_to_bit_it_10_vnu_83_in_2, msg_to_bit_it_10_vnu_84_in_0, msg_to_bit_it_10_vnu_84_in_1, msg_to_bit_it_10_vnu_84_in_2, msg_to_bit_it_10_vnu_85_in_0, msg_to_bit_it_10_vnu_85_in_1, msg_to_bit_it_10_vnu_85_in_2, msg_to_bit_it_10_vnu_86_in_0, msg_to_bit_it_10_vnu_86_in_1, msg_to_bit_it_10_vnu_86_in_2, msg_to_bit_it_10_vnu_87_in_0, msg_to_bit_it_10_vnu_87_in_1, msg_to_bit_it_10_vnu_87_in_2, msg_to_bit_it_10_vnu_88_in_0, msg_to_bit_it_10_vnu_88_in_1, msg_to_bit_it_10_vnu_88_in_2, msg_to_bit_it_10_vnu_89_in_0, msg_to_bit_it_10_vnu_89_in_1, msg_to_bit_it_10_vnu_89_in_2, msg_to_bit_it_10_vnu_90_in_0, msg_to_bit_it_10_vnu_90_in_1, msg_to_bit_it_10_vnu_90_in_2, msg_to_bit_it_10_vnu_91_in_0, msg_to_bit_it_10_vnu_91_in_1, msg_to_bit_it_10_vnu_91_in_2, msg_to_bit_it_10_vnu_92_in_0, msg_to_bit_it_10_vnu_92_in_1, msg_to_bit_it_10_vnu_92_in_2, msg_to_bit_it_10_vnu_93_in_0, msg_to_bit_it_10_vnu_93_in_1, msg_to_bit_it_10_vnu_93_in_2, msg_to_bit_it_10_vnu_94_in_0, msg_to_bit_it_10_vnu_94_in_1, msg_to_bit_it_10_vnu_94_in_2, msg_to_bit_it_10_vnu_95_in_0, msg_to_bit_it_10_vnu_95_in_1, msg_to_bit_it_10_vnu_95_in_2, msg_to_bit_it_10_vnu_96_in_0, msg_to_bit_it_10_vnu_96_in_1, msg_to_bit_it_10_vnu_96_in_2, msg_to_bit_it_10_vnu_97_in_0, msg_to_bit_it_10_vnu_97_in_1, msg_to_bit_it_10_vnu_97_in_2, msg_to_bit_it_10_vnu_98_in_0, msg_to_bit_it_10_vnu_98_in_1, msg_to_bit_it_10_vnu_98_in_2, msg_to_bit_it_10_vnu_99_in_0, msg_to_bit_it_10_vnu_99_in_1, msg_to_bit_it_10_vnu_99_in_2, msg_to_bit_it_10_vnu_100_in_0, msg_to_bit_it_10_vnu_100_in_1, msg_to_bit_it_10_vnu_100_in_2, msg_to_bit_it_10_vnu_101_in_0, msg_to_bit_it_10_vnu_101_in_1, msg_to_bit_it_10_vnu_101_in_2, msg_to_bit_it_10_vnu_102_in_0, msg_to_bit_it_10_vnu_102_in_1, msg_to_bit_it_10_vnu_102_in_2, msg_to_bit_it_10_vnu_103_in_0, msg_to_bit_it_10_vnu_103_in_1, msg_to_bit_it_10_vnu_103_in_2, msg_to_bit_it_10_vnu_104_in_0, msg_to_bit_it_10_vnu_104_in_1, msg_to_bit_it_10_vnu_104_in_2, msg_to_bit_it_10_vnu_105_in_0, msg_to_bit_it_10_vnu_105_in_1, msg_to_bit_it_10_vnu_105_in_2, msg_to_bit_it_10_vnu_106_in_0, msg_to_bit_it_10_vnu_106_in_1, msg_to_bit_it_10_vnu_106_in_2, msg_to_bit_it_10_vnu_107_in_0, msg_to_bit_it_10_vnu_107_in_1, msg_to_bit_it_10_vnu_107_in_2, msg_to_bit_it_10_vnu_108_in_0, msg_to_bit_it_10_vnu_108_in_1, msg_to_bit_it_10_vnu_108_in_2, msg_to_bit_it_10_vnu_109_in_0, msg_to_bit_it_10_vnu_109_in_1, msg_to_bit_it_10_vnu_109_in_2, msg_to_bit_it_10_vnu_110_in_0, msg_to_bit_it_10_vnu_110_in_1, msg_to_bit_it_10_vnu_110_in_2, msg_to_bit_it_10_vnu_111_in_0, msg_to_bit_it_10_vnu_111_in_1, msg_to_bit_it_10_vnu_111_in_2, msg_to_bit_it_10_vnu_112_in_0, msg_to_bit_it_10_vnu_112_in_1, msg_to_bit_it_10_vnu_112_in_2, msg_to_bit_it_10_vnu_113_in_0, msg_to_bit_it_10_vnu_113_in_1, msg_to_bit_it_10_vnu_113_in_2, msg_to_bit_it_10_vnu_114_in_0, msg_to_bit_it_10_vnu_114_in_1, msg_to_bit_it_10_vnu_114_in_2, msg_to_bit_it_10_vnu_115_in_0, msg_to_bit_it_10_vnu_115_in_1, msg_to_bit_it_10_vnu_115_in_2, msg_to_bit_it_10_vnu_116_in_0, msg_to_bit_it_10_vnu_116_in_1, msg_to_bit_it_10_vnu_116_in_2, msg_to_bit_it_10_vnu_117_in_0, msg_to_bit_it_10_vnu_117_in_1, msg_to_bit_it_10_vnu_117_in_2, msg_to_bit_it_10_vnu_118_in_0, msg_to_bit_it_10_vnu_118_in_1, msg_to_bit_it_10_vnu_118_in_2, msg_to_bit_it_10_vnu_119_in_0, msg_to_bit_it_10_vnu_119_in_1, msg_to_bit_it_10_vnu_119_in_2, msg_to_bit_it_10_vnu_120_in_0, msg_to_bit_it_10_vnu_120_in_1, msg_to_bit_it_10_vnu_120_in_2, msg_to_bit_it_10_vnu_121_in_0, msg_to_bit_it_10_vnu_121_in_1, msg_to_bit_it_10_vnu_121_in_2, msg_to_bit_it_10_vnu_122_in_0, msg_to_bit_it_10_vnu_122_in_1, msg_to_bit_it_10_vnu_122_in_2, msg_to_bit_it_10_vnu_123_in_0, msg_to_bit_it_10_vnu_123_in_1, msg_to_bit_it_10_vnu_123_in_2, msg_to_bit_it_10_vnu_124_in_0, msg_to_bit_it_10_vnu_124_in_1, msg_to_bit_it_10_vnu_124_in_2, msg_to_bit_it_10_vnu_125_in_0, msg_to_bit_it_10_vnu_125_in_1, msg_to_bit_it_10_vnu_125_in_2, msg_to_bit_it_10_vnu_126_in_0, msg_to_bit_it_10_vnu_126_in_1, msg_to_bit_it_10_vnu_126_in_2, msg_to_bit_it_10_vnu_127_in_0, msg_to_bit_it_10_vnu_127_in_1, msg_to_bit_it_10_vnu_127_in_2, msg_to_bit_it_10_vnu_128_in_0, msg_to_bit_it_10_vnu_128_in_1, msg_to_bit_it_10_vnu_128_in_2, msg_to_bit_it_10_vnu_129_in_0, msg_to_bit_it_10_vnu_129_in_1, msg_to_bit_it_10_vnu_129_in_2, msg_to_bit_it_10_vnu_130_in_0, msg_to_bit_it_10_vnu_130_in_1, msg_to_bit_it_10_vnu_130_in_2, msg_to_bit_it_10_vnu_131_in_0, msg_to_bit_it_10_vnu_131_in_1, msg_to_bit_it_10_vnu_131_in_2, msg_to_bit_it_10_vnu_132_in_0, msg_to_bit_it_10_vnu_132_in_1, msg_to_bit_it_10_vnu_132_in_2, msg_to_bit_it_10_vnu_133_in_0, msg_to_bit_it_10_vnu_133_in_1, msg_to_bit_it_10_vnu_133_in_2, msg_to_bit_it_10_vnu_134_in_0, msg_to_bit_it_10_vnu_134_in_1, msg_to_bit_it_10_vnu_134_in_2, msg_to_bit_it_10_vnu_135_in_0, msg_to_bit_it_10_vnu_135_in_1, msg_to_bit_it_10_vnu_135_in_2, msg_to_bit_it_10_vnu_136_in_0, msg_to_bit_it_10_vnu_136_in_1, msg_to_bit_it_10_vnu_136_in_2, msg_to_bit_it_10_vnu_137_in_0, msg_to_bit_it_10_vnu_137_in_1, msg_to_bit_it_10_vnu_137_in_2, msg_to_bit_it_10_vnu_138_in_0, msg_to_bit_it_10_vnu_138_in_1, msg_to_bit_it_10_vnu_138_in_2, msg_to_bit_it_10_vnu_139_in_0, msg_to_bit_it_10_vnu_139_in_1, msg_to_bit_it_10_vnu_139_in_2, msg_to_bit_it_10_vnu_140_in_0, msg_to_bit_it_10_vnu_140_in_1, msg_to_bit_it_10_vnu_140_in_2, msg_to_bit_it_10_vnu_141_in_0, msg_to_bit_it_10_vnu_141_in_1, msg_to_bit_it_10_vnu_141_in_2, msg_to_bit_it_10_vnu_142_in_0, msg_to_bit_it_10_vnu_142_in_1, msg_to_bit_it_10_vnu_142_in_2, msg_to_bit_it_10_vnu_143_in_0, msg_to_bit_it_10_vnu_143_in_1, msg_to_bit_it_10_vnu_143_in_2, msg_to_bit_it_10_vnu_144_in_0, msg_to_bit_it_10_vnu_144_in_1, msg_to_bit_it_10_vnu_144_in_2, msg_to_bit_it_10_vnu_145_in_0, msg_to_bit_it_10_vnu_145_in_1, msg_to_bit_it_10_vnu_145_in_2, msg_to_bit_it_10_vnu_146_in_0, msg_to_bit_it_10_vnu_146_in_1, msg_to_bit_it_10_vnu_146_in_2, msg_to_bit_it_10_vnu_147_in_0, msg_to_bit_it_10_vnu_147_in_1, msg_to_bit_it_10_vnu_147_in_2, msg_to_bit_it_10_vnu_148_in_0, msg_to_bit_it_10_vnu_148_in_1, msg_to_bit_it_10_vnu_148_in_2, msg_to_bit_it_10_vnu_149_in_0, msg_to_bit_it_10_vnu_149_in_1, msg_to_bit_it_10_vnu_149_in_2, msg_to_bit_it_10_vnu_150_in_0, msg_to_bit_it_10_vnu_150_in_1, msg_to_bit_it_10_vnu_150_in_2, msg_to_bit_it_10_vnu_151_in_0, msg_to_bit_it_10_vnu_151_in_1, msg_to_bit_it_10_vnu_151_in_2, msg_to_bit_it_10_vnu_152_in_0, msg_to_bit_it_10_vnu_152_in_1, msg_to_bit_it_10_vnu_152_in_2, msg_to_bit_it_10_vnu_153_in_0, msg_to_bit_it_10_vnu_153_in_1, msg_to_bit_it_10_vnu_153_in_2, msg_to_bit_it_10_vnu_154_in_0, msg_to_bit_it_10_vnu_154_in_1, msg_to_bit_it_10_vnu_154_in_2, msg_to_bit_it_10_vnu_155_in_0, msg_to_bit_it_10_vnu_155_in_1, msg_to_bit_it_10_vnu_155_in_2, msg_to_bit_it_10_vnu_156_in_0, msg_to_bit_it_10_vnu_156_in_1, msg_to_bit_it_10_vnu_156_in_2, msg_to_bit_it_10_vnu_157_in_0, msg_to_bit_it_10_vnu_157_in_1, msg_to_bit_it_10_vnu_157_in_2, msg_to_bit_it_10_vnu_158_in_0, msg_to_bit_it_10_vnu_158_in_1, msg_to_bit_it_10_vnu_158_in_2, msg_to_bit_it_10_vnu_159_in_0, msg_to_bit_it_10_vnu_159_in_1, msg_to_bit_it_10_vnu_159_in_2, msg_to_bit_it_10_vnu_160_in_0, msg_to_bit_it_10_vnu_160_in_1, msg_to_bit_it_10_vnu_160_in_2, msg_to_bit_it_10_vnu_161_in_0, msg_to_bit_it_10_vnu_161_in_1, msg_to_bit_it_10_vnu_161_in_2, msg_to_bit_it_10_vnu_162_in_0, msg_to_bit_it_10_vnu_162_in_1, msg_to_bit_it_10_vnu_162_in_2, msg_to_bit_it_10_vnu_163_in_0, msg_to_bit_it_10_vnu_163_in_1, msg_to_bit_it_10_vnu_163_in_2, msg_to_bit_it_10_vnu_164_in_0, msg_to_bit_it_10_vnu_164_in_1, msg_to_bit_it_10_vnu_164_in_2, msg_to_bit_it_10_vnu_165_in_0, msg_to_bit_it_10_vnu_165_in_1, msg_to_bit_it_10_vnu_165_in_2, msg_to_bit_it_10_vnu_166_in_0, msg_to_bit_it_10_vnu_166_in_1, msg_to_bit_it_10_vnu_166_in_2, msg_to_bit_it_10_vnu_167_in_0, msg_to_bit_it_10_vnu_167_in_1, msg_to_bit_it_10_vnu_167_in_2, msg_to_bit_it_10_vnu_168_in_0, msg_to_bit_it_10_vnu_168_in_1, msg_to_bit_it_10_vnu_168_in_2, msg_to_bit_it_10_vnu_169_in_0, msg_to_bit_it_10_vnu_169_in_1, msg_to_bit_it_10_vnu_169_in_2, msg_to_bit_it_10_vnu_170_in_0, msg_to_bit_it_10_vnu_170_in_1, msg_to_bit_it_10_vnu_170_in_2, msg_to_bit_it_10_vnu_171_in_0, msg_to_bit_it_10_vnu_171_in_1, msg_to_bit_it_10_vnu_171_in_2, msg_to_bit_it_10_vnu_172_in_0, msg_to_bit_it_10_vnu_172_in_1, msg_to_bit_it_10_vnu_172_in_2, msg_to_bit_it_10_vnu_173_in_0, msg_to_bit_it_10_vnu_173_in_1, msg_to_bit_it_10_vnu_173_in_2, msg_to_bit_it_10_vnu_174_in_0, msg_to_bit_it_10_vnu_174_in_1, msg_to_bit_it_10_vnu_174_in_2, msg_to_bit_it_10_vnu_175_in_0, msg_to_bit_it_10_vnu_175_in_1, msg_to_bit_it_10_vnu_175_in_2, msg_to_bit_it_10_vnu_176_in_0, msg_to_bit_it_10_vnu_176_in_1, msg_to_bit_it_10_vnu_176_in_2, msg_to_bit_it_10_vnu_177_in_0, msg_to_bit_it_10_vnu_177_in_1, msg_to_bit_it_10_vnu_177_in_2, msg_to_bit_it_10_vnu_178_in_0, msg_to_bit_it_10_vnu_178_in_1, msg_to_bit_it_10_vnu_178_in_2, msg_to_bit_it_10_vnu_179_in_0, msg_to_bit_it_10_vnu_179_in_1, msg_to_bit_it_10_vnu_179_in_2, msg_to_bit_it_10_vnu_180_in_0, msg_to_bit_it_10_vnu_180_in_1, msg_to_bit_it_10_vnu_180_in_2, msg_to_bit_it_10_vnu_181_in_0, msg_to_bit_it_10_vnu_181_in_1, msg_to_bit_it_10_vnu_181_in_2, msg_to_bit_it_10_vnu_182_in_0, msg_to_bit_it_10_vnu_182_in_1, msg_to_bit_it_10_vnu_182_in_2, msg_to_bit_it_10_vnu_183_in_0, msg_to_bit_it_10_vnu_183_in_1, msg_to_bit_it_10_vnu_183_in_2, msg_to_bit_it_10_vnu_184_in_0, msg_to_bit_it_10_vnu_184_in_1, msg_to_bit_it_10_vnu_184_in_2, msg_to_bit_it_10_vnu_185_in_0, msg_to_bit_it_10_vnu_185_in_1, msg_to_bit_it_10_vnu_185_in_2, msg_to_bit_it_10_vnu_186_in_0, msg_to_bit_it_10_vnu_186_in_1, msg_to_bit_it_10_vnu_186_in_2, msg_to_bit_it_10_vnu_187_in_0, msg_to_bit_it_10_vnu_187_in_1, msg_to_bit_it_10_vnu_187_in_2, msg_to_bit_it_10_vnu_188_in_0, msg_to_bit_it_10_vnu_188_in_1, msg_to_bit_it_10_vnu_188_in_2, msg_to_bit_it_10_vnu_189_in_0, msg_to_bit_it_10_vnu_189_in_1, msg_to_bit_it_10_vnu_189_in_2, msg_to_bit_it_10_vnu_190_in_0, msg_to_bit_it_10_vnu_190_in_1, msg_to_bit_it_10_vnu_190_in_2, msg_to_bit_it_10_vnu_191_in_0, msg_to_bit_it_10_vnu_191_in_1, msg_to_bit_it_10_vnu_191_in_2, msg_to_bit_it_10_vnu_192_in_0, msg_to_bit_it_10_vnu_192_in_1, msg_to_bit_it_10_vnu_192_in_2, msg_to_bit_it_10_vnu_193_in_0, msg_to_bit_it_10_vnu_193_in_1, msg_to_bit_it_10_vnu_193_in_2, msg_to_bit_it_10_vnu_194_in_0, msg_to_bit_it_10_vnu_194_in_1, msg_to_bit_it_10_vnu_194_in_2, msg_to_bit_it_10_vnu_195_in_0, msg_to_bit_it_10_vnu_195_in_1, msg_to_bit_it_10_vnu_195_in_2, msg_to_bit_it_10_vnu_196_in_0, msg_to_bit_it_10_vnu_196_in_1, msg_to_bit_it_10_vnu_196_in_2, msg_to_bit_it_10_vnu_197_in_0, msg_to_bit_it_10_vnu_197_in_1, msg_to_bit_it_10_vnu_197_in_2, msg_to_bit_it_11_vnu_0_in_0, msg_to_bit_it_11_vnu_0_in_1, msg_to_bit_it_11_vnu_0_in_2, msg_to_bit_it_11_vnu_1_in_0, msg_to_bit_it_11_vnu_1_in_1, msg_to_bit_it_11_vnu_1_in_2, msg_to_bit_it_11_vnu_2_in_0, msg_to_bit_it_11_vnu_2_in_1, msg_to_bit_it_11_vnu_2_in_2, msg_to_bit_it_11_vnu_3_in_0, msg_to_bit_it_11_vnu_3_in_1, msg_to_bit_it_11_vnu_3_in_2, msg_to_bit_it_11_vnu_4_in_0, msg_to_bit_it_11_vnu_4_in_1, msg_to_bit_it_11_vnu_4_in_2, msg_to_bit_it_11_vnu_5_in_0, msg_to_bit_it_11_vnu_5_in_1, msg_to_bit_it_11_vnu_5_in_2, msg_to_bit_it_11_vnu_6_in_0, msg_to_bit_it_11_vnu_6_in_1, msg_to_bit_it_11_vnu_6_in_2, msg_to_bit_it_11_vnu_7_in_0, msg_to_bit_it_11_vnu_7_in_1, msg_to_bit_it_11_vnu_7_in_2, msg_to_bit_it_11_vnu_8_in_0, msg_to_bit_it_11_vnu_8_in_1, msg_to_bit_it_11_vnu_8_in_2, msg_to_bit_it_11_vnu_9_in_0, msg_to_bit_it_11_vnu_9_in_1, msg_to_bit_it_11_vnu_9_in_2, msg_to_bit_it_11_vnu_10_in_0, msg_to_bit_it_11_vnu_10_in_1, msg_to_bit_it_11_vnu_10_in_2, msg_to_bit_it_11_vnu_11_in_0, msg_to_bit_it_11_vnu_11_in_1, msg_to_bit_it_11_vnu_11_in_2, msg_to_bit_it_11_vnu_12_in_0, msg_to_bit_it_11_vnu_12_in_1, msg_to_bit_it_11_vnu_12_in_2, msg_to_bit_it_11_vnu_13_in_0, msg_to_bit_it_11_vnu_13_in_1, msg_to_bit_it_11_vnu_13_in_2, msg_to_bit_it_11_vnu_14_in_0, msg_to_bit_it_11_vnu_14_in_1, msg_to_bit_it_11_vnu_14_in_2, msg_to_bit_it_11_vnu_15_in_0, msg_to_bit_it_11_vnu_15_in_1, msg_to_bit_it_11_vnu_15_in_2, msg_to_bit_it_11_vnu_16_in_0, msg_to_bit_it_11_vnu_16_in_1, msg_to_bit_it_11_vnu_16_in_2, msg_to_bit_it_11_vnu_17_in_0, msg_to_bit_it_11_vnu_17_in_1, msg_to_bit_it_11_vnu_17_in_2, msg_to_bit_it_11_vnu_18_in_0, msg_to_bit_it_11_vnu_18_in_1, msg_to_bit_it_11_vnu_18_in_2, msg_to_bit_it_11_vnu_19_in_0, msg_to_bit_it_11_vnu_19_in_1, msg_to_bit_it_11_vnu_19_in_2, msg_to_bit_it_11_vnu_20_in_0, msg_to_bit_it_11_vnu_20_in_1, msg_to_bit_it_11_vnu_20_in_2, msg_to_bit_it_11_vnu_21_in_0, msg_to_bit_it_11_vnu_21_in_1, msg_to_bit_it_11_vnu_21_in_2, msg_to_bit_it_11_vnu_22_in_0, msg_to_bit_it_11_vnu_22_in_1, msg_to_bit_it_11_vnu_22_in_2, msg_to_bit_it_11_vnu_23_in_0, msg_to_bit_it_11_vnu_23_in_1, msg_to_bit_it_11_vnu_23_in_2, msg_to_bit_it_11_vnu_24_in_0, msg_to_bit_it_11_vnu_24_in_1, msg_to_bit_it_11_vnu_24_in_2, msg_to_bit_it_11_vnu_25_in_0, msg_to_bit_it_11_vnu_25_in_1, msg_to_bit_it_11_vnu_25_in_2, msg_to_bit_it_11_vnu_26_in_0, msg_to_bit_it_11_vnu_26_in_1, msg_to_bit_it_11_vnu_26_in_2, msg_to_bit_it_11_vnu_27_in_0, msg_to_bit_it_11_vnu_27_in_1, msg_to_bit_it_11_vnu_27_in_2, msg_to_bit_it_11_vnu_28_in_0, msg_to_bit_it_11_vnu_28_in_1, msg_to_bit_it_11_vnu_28_in_2, msg_to_bit_it_11_vnu_29_in_0, msg_to_bit_it_11_vnu_29_in_1, msg_to_bit_it_11_vnu_29_in_2, msg_to_bit_it_11_vnu_30_in_0, msg_to_bit_it_11_vnu_30_in_1, msg_to_bit_it_11_vnu_30_in_2, msg_to_bit_it_11_vnu_31_in_0, msg_to_bit_it_11_vnu_31_in_1, msg_to_bit_it_11_vnu_31_in_2, msg_to_bit_it_11_vnu_32_in_0, msg_to_bit_it_11_vnu_32_in_1, msg_to_bit_it_11_vnu_32_in_2, msg_to_bit_it_11_vnu_33_in_0, msg_to_bit_it_11_vnu_33_in_1, msg_to_bit_it_11_vnu_33_in_2, msg_to_bit_it_11_vnu_34_in_0, msg_to_bit_it_11_vnu_34_in_1, msg_to_bit_it_11_vnu_34_in_2, msg_to_bit_it_11_vnu_35_in_0, msg_to_bit_it_11_vnu_35_in_1, msg_to_bit_it_11_vnu_35_in_2, msg_to_bit_it_11_vnu_36_in_0, msg_to_bit_it_11_vnu_36_in_1, msg_to_bit_it_11_vnu_36_in_2, msg_to_bit_it_11_vnu_37_in_0, msg_to_bit_it_11_vnu_37_in_1, msg_to_bit_it_11_vnu_37_in_2, msg_to_bit_it_11_vnu_38_in_0, msg_to_bit_it_11_vnu_38_in_1, msg_to_bit_it_11_vnu_38_in_2, msg_to_bit_it_11_vnu_39_in_0, msg_to_bit_it_11_vnu_39_in_1, msg_to_bit_it_11_vnu_39_in_2, msg_to_bit_it_11_vnu_40_in_0, msg_to_bit_it_11_vnu_40_in_1, msg_to_bit_it_11_vnu_40_in_2, msg_to_bit_it_11_vnu_41_in_0, msg_to_bit_it_11_vnu_41_in_1, msg_to_bit_it_11_vnu_41_in_2, msg_to_bit_it_11_vnu_42_in_0, msg_to_bit_it_11_vnu_42_in_1, msg_to_bit_it_11_vnu_42_in_2, msg_to_bit_it_11_vnu_43_in_0, msg_to_bit_it_11_vnu_43_in_1, msg_to_bit_it_11_vnu_43_in_2, msg_to_bit_it_11_vnu_44_in_0, msg_to_bit_it_11_vnu_44_in_1, msg_to_bit_it_11_vnu_44_in_2, msg_to_bit_it_11_vnu_45_in_0, msg_to_bit_it_11_vnu_45_in_1, msg_to_bit_it_11_vnu_45_in_2, msg_to_bit_it_11_vnu_46_in_0, msg_to_bit_it_11_vnu_46_in_1, msg_to_bit_it_11_vnu_46_in_2, msg_to_bit_it_11_vnu_47_in_0, msg_to_bit_it_11_vnu_47_in_1, msg_to_bit_it_11_vnu_47_in_2, msg_to_bit_it_11_vnu_48_in_0, msg_to_bit_it_11_vnu_48_in_1, msg_to_bit_it_11_vnu_48_in_2, msg_to_bit_it_11_vnu_49_in_0, msg_to_bit_it_11_vnu_49_in_1, msg_to_bit_it_11_vnu_49_in_2, msg_to_bit_it_11_vnu_50_in_0, msg_to_bit_it_11_vnu_50_in_1, msg_to_bit_it_11_vnu_50_in_2, msg_to_bit_it_11_vnu_51_in_0, msg_to_bit_it_11_vnu_51_in_1, msg_to_bit_it_11_vnu_51_in_2, msg_to_bit_it_11_vnu_52_in_0, msg_to_bit_it_11_vnu_52_in_1, msg_to_bit_it_11_vnu_52_in_2, msg_to_bit_it_11_vnu_53_in_0, msg_to_bit_it_11_vnu_53_in_1, msg_to_bit_it_11_vnu_53_in_2, msg_to_bit_it_11_vnu_54_in_0, msg_to_bit_it_11_vnu_54_in_1, msg_to_bit_it_11_vnu_54_in_2, msg_to_bit_it_11_vnu_55_in_0, msg_to_bit_it_11_vnu_55_in_1, msg_to_bit_it_11_vnu_55_in_2, msg_to_bit_it_11_vnu_56_in_0, msg_to_bit_it_11_vnu_56_in_1, msg_to_bit_it_11_vnu_56_in_2, msg_to_bit_it_11_vnu_57_in_0, msg_to_bit_it_11_vnu_57_in_1, msg_to_bit_it_11_vnu_57_in_2, msg_to_bit_it_11_vnu_58_in_0, msg_to_bit_it_11_vnu_58_in_1, msg_to_bit_it_11_vnu_58_in_2, msg_to_bit_it_11_vnu_59_in_0, msg_to_bit_it_11_vnu_59_in_1, msg_to_bit_it_11_vnu_59_in_2, msg_to_bit_it_11_vnu_60_in_0, msg_to_bit_it_11_vnu_60_in_1, msg_to_bit_it_11_vnu_60_in_2, msg_to_bit_it_11_vnu_61_in_0, msg_to_bit_it_11_vnu_61_in_1, msg_to_bit_it_11_vnu_61_in_2, msg_to_bit_it_11_vnu_62_in_0, msg_to_bit_it_11_vnu_62_in_1, msg_to_bit_it_11_vnu_62_in_2, msg_to_bit_it_11_vnu_63_in_0, msg_to_bit_it_11_vnu_63_in_1, msg_to_bit_it_11_vnu_63_in_2, msg_to_bit_it_11_vnu_64_in_0, msg_to_bit_it_11_vnu_64_in_1, msg_to_bit_it_11_vnu_64_in_2, msg_to_bit_it_11_vnu_65_in_0, msg_to_bit_it_11_vnu_65_in_1, msg_to_bit_it_11_vnu_65_in_2, msg_to_bit_it_11_vnu_66_in_0, msg_to_bit_it_11_vnu_66_in_1, msg_to_bit_it_11_vnu_66_in_2, msg_to_bit_it_11_vnu_67_in_0, msg_to_bit_it_11_vnu_67_in_1, msg_to_bit_it_11_vnu_67_in_2, msg_to_bit_it_11_vnu_68_in_0, msg_to_bit_it_11_vnu_68_in_1, msg_to_bit_it_11_vnu_68_in_2, msg_to_bit_it_11_vnu_69_in_0, msg_to_bit_it_11_vnu_69_in_1, msg_to_bit_it_11_vnu_69_in_2, msg_to_bit_it_11_vnu_70_in_0, msg_to_bit_it_11_vnu_70_in_1, msg_to_bit_it_11_vnu_70_in_2, msg_to_bit_it_11_vnu_71_in_0, msg_to_bit_it_11_vnu_71_in_1, msg_to_bit_it_11_vnu_71_in_2, msg_to_bit_it_11_vnu_72_in_0, msg_to_bit_it_11_vnu_72_in_1, msg_to_bit_it_11_vnu_72_in_2, msg_to_bit_it_11_vnu_73_in_0, msg_to_bit_it_11_vnu_73_in_1, msg_to_bit_it_11_vnu_73_in_2, msg_to_bit_it_11_vnu_74_in_0, msg_to_bit_it_11_vnu_74_in_1, msg_to_bit_it_11_vnu_74_in_2, msg_to_bit_it_11_vnu_75_in_0, msg_to_bit_it_11_vnu_75_in_1, msg_to_bit_it_11_vnu_75_in_2, msg_to_bit_it_11_vnu_76_in_0, msg_to_bit_it_11_vnu_76_in_1, msg_to_bit_it_11_vnu_76_in_2, msg_to_bit_it_11_vnu_77_in_0, msg_to_bit_it_11_vnu_77_in_1, msg_to_bit_it_11_vnu_77_in_2, msg_to_bit_it_11_vnu_78_in_0, msg_to_bit_it_11_vnu_78_in_1, msg_to_bit_it_11_vnu_78_in_2, msg_to_bit_it_11_vnu_79_in_0, msg_to_bit_it_11_vnu_79_in_1, msg_to_bit_it_11_vnu_79_in_2, msg_to_bit_it_11_vnu_80_in_0, msg_to_bit_it_11_vnu_80_in_1, msg_to_bit_it_11_vnu_80_in_2, msg_to_bit_it_11_vnu_81_in_0, msg_to_bit_it_11_vnu_81_in_1, msg_to_bit_it_11_vnu_81_in_2, msg_to_bit_it_11_vnu_82_in_0, msg_to_bit_it_11_vnu_82_in_1, msg_to_bit_it_11_vnu_82_in_2, msg_to_bit_it_11_vnu_83_in_0, msg_to_bit_it_11_vnu_83_in_1, msg_to_bit_it_11_vnu_83_in_2, msg_to_bit_it_11_vnu_84_in_0, msg_to_bit_it_11_vnu_84_in_1, msg_to_bit_it_11_vnu_84_in_2, msg_to_bit_it_11_vnu_85_in_0, msg_to_bit_it_11_vnu_85_in_1, msg_to_bit_it_11_vnu_85_in_2, msg_to_bit_it_11_vnu_86_in_0, msg_to_bit_it_11_vnu_86_in_1, msg_to_bit_it_11_vnu_86_in_2, msg_to_bit_it_11_vnu_87_in_0, msg_to_bit_it_11_vnu_87_in_1, msg_to_bit_it_11_vnu_87_in_2, msg_to_bit_it_11_vnu_88_in_0, msg_to_bit_it_11_vnu_88_in_1, msg_to_bit_it_11_vnu_88_in_2, msg_to_bit_it_11_vnu_89_in_0, msg_to_bit_it_11_vnu_89_in_1, msg_to_bit_it_11_vnu_89_in_2, msg_to_bit_it_11_vnu_90_in_0, msg_to_bit_it_11_vnu_90_in_1, msg_to_bit_it_11_vnu_90_in_2, msg_to_bit_it_11_vnu_91_in_0, msg_to_bit_it_11_vnu_91_in_1, msg_to_bit_it_11_vnu_91_in_2, msg_to_bit_it_11_vnu_92_in_0, msg_to_bit_it_11_vnu_92_in_1, msg_to_bit_it_11_vnu_92_in_2, msg_to_bit_it_11_vnu_93_in_0, msg_to_bit_it_11_vnu_93_in_1, msg_to_bit_it_11_vnu_93_in_2, msg_to_bit_it_11_vnu_94_in_0, msg_to_bit_it_11_vnu_94_in_1, msg_to_bit_it_11_vnu_94_in_2, msg_to_bit_it_11_vnu_95_in_0, msg_to_bit_it_11_vnu_95_in_1, msg_to_bit_it_11_vnu_95_in_2, msg_to_bit_it_11_vnu_96_in_0, msg_to_bit_it_11_vnu_96_in_1, msg_to_bit_it_11_vnu_96_in_2, msg_to_bit_it_11_vnu_97_in_0, msg_to_bit_it_11_vnu_97_in_1, msg_to_bit_it_11_vnu_97_in_2, msg_to_bit_it_11_vnu_98_in_0, msg_to_bit_it_11_vnu_98_in_1, msg_to_bit_it_11_vnu_98_in_2, msg_to_bit_it_11_vnu_99_in_0, msg_to_bit_it_11_vnu_99_in_1, msg_to_bit_it_11_vnu_99_in_2, msg_to_bit_it_11_vnu_100_in_0, msg_to_bit_it_11_vnu_100_in_1, msg_to_bit_it_11_vnu_100_in_2, msg_to_bit_it_11_vnu_101_in_0, msg_to_bit_it_11_vnu_101_in_1, msg_to_bit_it_11_vnu_101_in_2, msg_to_bit_it_11_vnu_102_in_0, msg_to_bit_it_11_vnu_102_in_1, msg_to_bit_it_11_vnu_102_in_2, msg_to_bit_it_11_vnu_103_in_0, msg_to_bit_it_11_vnu_103_in_1, msg_to_bit_it_11_vnu_103_in_2, msg_to_bit_it_11_vnu_104_in_0, msg_to_bit_it_11_vnu_104_in_1, msg_to_bit_it_11_vnu_104_in_2, msg_to_bit_it_11_vnu_105_in_0, msg_to_bit_it_11_vnu_105_in_1, msg_to_bit_it_11_vnu_105_in_2, msg_to_bit_it_11_vnu_106_in_0, msg_to_bit_it_11_vnu_106_in_1, msg_to_bit_it_11_vnu_106_in_2, msg_to_bit_it_11_vnu_107_in_0, msg_to_bit_it_11_vnu_107_in_1, msg_to_bit_it_11_vnu_107_in_2, msg_to_bit_it_11_vnu_108_in_0, msg_to_bit_it_11_vnu_108_in_1, msg_to_bit_it_11_vnu_108_in_2, msg_to_bit_it_11_vnu_109_in_0, msg_to_bit_it_11_vnu_109_in_1, msg_to_bit_it_11_vnu_109_in_2, msg_to_bit_it_11_vnu_110_in_0, msg_to_bit_it_11_vnu_110_in_1, msg_to_bit_it_11_vnu_110_in_2, msg_to_bit_it_11_vnu_111_in_0, msg_to_bit_it_11_vnu_111_in_1, msg_to_bit_it_11_vnu_111_in_2, msg_to_bit_it_11_vnu_112_in_0, msg_to_bit_it_11_vnu_112_in_1, msg_to_bit_it_11_vnu_112_in_2, msg_to_bit_it_11_vnu_113_in_0, msg_to_bit_it_11_vnu_113_in_1, msg_to_bit_it_11_vnu_113_in_2, msg_to_bit_it_11_vnu_114_in_0, msg_to_bit_it_11_vnu_114_in_1, msg_to_bit_it_11_vnu_114_in_2, msg_to_bit_it_11_vnu_115_in_0, msg_to_bit_it_11_vnu_115_in_1, msg_to_bit_it_11_vnu_115_in_2, msg_to_bit_it_11_vnu_116_in_0, msg_to_bit_it_11_vnu_116_in_1, msg_to_bit_it_11_vnu_116_in_2, msg_to_bit_it_11_vnu_117_in_0, msg_to_bit_it_11_vnu_117_in_1, msg_to_bit_it_11_vnu_117_in_2, msg_to_bit_it_11_vnu_118_in_0, msg_to_bit_it_11_vnu_118_in_1, msg_to_bit_it_11_vnu_118_in_2, msg_to_bit_it_11_vnu_119_in_0, msg_to_bit_it_11_vnu_119_in_1, msg_to_bit_it_11_vnu_119_in_2, msg_to_bit_it_11_vnu_120_in_0, msg_to_bit_it_11_vnu_120_in_1, msg_to_bit_it_11_vnu_120_in_2, msg_to_bit_it_11_vnu_121_in_0, msg_to_bit_it_11_vnu_121_in_1, msg_to_bit_it_11_vnu_121_in_2, msg_to_bit_it_11_vnu_122_in_0, msg_to_bit_it_11_vnu_122_in_1, msg_to_bit_it_11_vnu_122_in_2, msg_to_bit_it_11_vnu_123_in_0, msg_to_bit_it_11_vnu_123_in_1, msg_to_bit_it_11_vnu_123_in_2, msg_to_bit_it_11_vnu_124_in_0, msg_to_bit_it_11_vnu_124_in_1, msg_to_bit_it_11_vnu_124_in_2, msg_to_bit_it_11_vnu_125_in_0, msg_to_bit_it_11_vnu_125_in_1, msg_to_bit_it_11_vnu_125_in_2, msg_to_bit_it_11_vnu_126_in_0, msg_to_bit_it_11_vnu_126_in_1, msg_to_bit_it_11_vnu_126_in_2, msg_to_bit_it_11_vnu_127_in_0, msg_to_bit_it_11_vnu_127_in_1, msg_to_bit_it_11_vnu_127_in_2, msg_to_bit_it_11_vnu_128_in_0, msg_to_bit_it_11_vnu_128_in_1, msg_to_bit_it_11_vnu_128_in_2, msg_to_bit_it_11_vnu_129_in_0, msg_to_bit_it_11_vnu_129_in_1, msg_to_bit_it_11_vnu_129_in_2, msg_to_bit_it_11_vnu_130_in_0, msg_to_bit_it_11_vnu_130_in_1, msg_to_bit_it_11_vnu_130_in_2, msg_to_bit_it_11_vnu_131_in_0, msg_to_bit_it_11_vnu_131_in_1, msg_to_bit_it_11_vnu_131_in_2, msg_to_bit_it_11_vnu_132_in_0, msg_to_bit_it_11_vnu_132_in_1, msg_to_bit_it_11_vnu_132_in_2, msg_to_bit_it_11_vnu_133_in_0, msg_to_bit_it_11_vnu_133_in_1, msg_to_bit_it_11_vnu_133_in_2, msg_to_bit_it_11_vnu_134_in_0, msg_to_bit_it_11_vnu_134_in_1, msg_to_bit_it_11_vnu_134_in_2, msg_to_bit_it_11_vnu_135_in_0, msg_to_bit_it_11_vnu_135_in_1, msg_to_bit_it_11_vnu_135_in_2, msg_to_bit_it_11_vnu_136_in_0, msg_to_bit_it_11_vnu_136_in_1, msg_to_bit_it_11_vnu_136_in_2, msg_to_bit_it_11_vnu_137_in_0, msg_to_bit_it_11_vnu_137_in_1, msg_to_bit_it_11_vnu_137_in_2, msg_to_bit_it_11_vnu_138_in_0, msg_to_bit_it_11_vnu_138_in_1, msg_to_bit_it_11_vnu_138_in_2, msg_to_bit_it_11_vnu_139_in_0, msg_to_bit_it_11_vnu_139_in_1, msg_to_bit_it_11_vnu_139_in_2, msg_to_bit_it_11_vnu_140_in_0, msg_to_bit_it_11_vnu_140_in_1, msg_to_bit_it_11_vnu_140_in_2, msg_to_bit_it_11_vnu_141_in_0, msg_to_bit_it_11_vnu_141_in_1, msg_to_bit_it_11_vnu_141_in_2, msg_to_bit_it_11_vnu_142_in_0, msg_to_bit_it_11_vnu_142_in_1, msg_to_bit_it_11_vnu_142_in_2, msg_to_bit_it_11_vnu_143_in_0, msg_to_bit_it_11_vnu_143_in_1, msg_to_bit_it_11_vnu_143_in_2, msg_to_bit_it_11_vnu_144_in_0, msg_to_bit_it_11_vnu_144_in_1, msg_to_bit_it_11_vnu_144_in_2, msg_to_bit_it_11_vnu_145_in_0, msg_to_bit_it_11_vnu_145_in_1, msg_to_bit_it_11_vnu_145_in_2, msg_to_bit_it_11_vnu_146_in_0, msg_to_bit_it_11_vnu_146_in_1, msg_to_bit_it_11_vnu_146_in_2, msg_to_bit_it_11_vnu_147_in_0, msg_to_bit_it_11_vnu_147_in_1, msg_to_bit_it_11_vnu_147_in_2, msg_to_bit_it_11_vnu_148_in_0, msg_to_bit_it_11_vnu_148_in_1, msg_to_bit_it_11_vnu_148_in_2, msg_to_bit_it_11_vnu_149_in_0, msg_to_bit_it_11_vnu_149_in_1, msg_to_bit_it_11_vnu_149_in_2, msg_to_bit_it_11_vnu_150_in_0, msg_to_bit_it_11_vnu_150_in_1, msg_to_bit_it_11_vnu_150_in_2, msg_to_bit_it_11_vnu_151_in_0, msg_to_bit_it_11_vnu_151_in_1, msg_to_bit_it_11_vnu_151_in_2, msg_to_bit_it_11_vnu_152_in_0, msg_to_bit_it_11_vnu_152_in_1, msg_to_bit_it_11_vnu_152_in_2, msg_to_bit_it_11_vnu_153_in_0, msg_to_bit_it_11_vnu_153_in_1, msg_to_bit_it_11_vnu_153_in_2, msg_to_bit_it_11_vnu_154_in_0, msg_to_bit_it_11_vnu_154_in_1, msg_to_bit_it_11_vnu_154_in_2, msg_to_bit_it_11_vnu_155_in_0, msg_to_bit_it_11_vnu_155_in_1, msg_to_bit_it_11_vnu_155_in_2, msg_to_bit_it_11_vnu_156_in_0, msg_to_bit_it_11_vnu_156_in_1, msg_to_bit_it_11_vnu_156_in_2, msg_to_bit_it_11_vnu_157_in_0, msg_to_bit_it_11_vnu_157_in_1, msg_to_bit_it_11_vnu_157_in_2, msg_to_bit_it_11_vnu_158_in_0, msg_to_bit_it_11_vnu_158_in_1, msg_to_bit_it_11_vnu_158_in_2, msg_to_bit_it_11_vnu_159_in_0, msg_to_bit_it_11_vnu_159_in_1, msg_to_bit_it_11_vnu_159_in_2, msg_to_bit_it_11_vnu_160_in_0, msg_to_bit_it_11_vnu_160_in_1, msg_to_bit_it_11_vnu_160_in_2, msg_to_bit_it_11_vnu_161_in_0, msg_to_bit_it_11_vnu_161_in_1, msg_to_bit_it_11_vnu_161_in_2, msg_to_bit_it_11_vnu_162_in_0, msg_to_bit_it_11_vnu_162_in_1, msg_to_bit_it_11_vnu_162_in_2, msg_to_bit_it_11_vnu_163_in_0, msg_to_bit_it_11_vnu_163_in_1, msg_to_bit_it_11_vnu_163_in_2, msg_to_bit_it_11_vnu_164_in_0, msg_to_bit_it_11_vnu_164_in_1, msg_to_bit_it_11_vnu_164_in_2, msg_to_bit_it_11_vnu_165_in_0, msg_to_bit_it_11_vnu_165_in_1, msg_to_bit_it_11_vnu_165_in_2, msg_to_bit_it_11_vnu_166_in_0, msg_to_bit_it_11_vnu_166_in_1, msg_to_bit_it_11_vnu_166_in_2, msg_to_bit_it_11_vnu_167_in_0, msg_to_bit_it_11_vnu_167_in_1, msg_to_bit_it_11_vnu_167_in_2, msg_to_bit_it_11_vnu_168_in_0, msg_to_bit_it_11_vnu_168_in_1, msg_to_bit_it_11_vnu_168_in_2, msg_to_bit_it_11_vnu_169_in_0, msg_to_bit_it_11_vnu_169_in_1, msg_to_bit_it_11_vnu_169_in_2, msg_to_bit_it_11_vnu_170_in_0, msg_to_bit_it_11_vnu_170_in_1, msg_to_bit_it_11_vnu_170_in_2, msg_to_bit_it_11_vnu_171_in_0, msg_to_bit_it_11_vnu_171_in_1, msg_to_bit_it_11_vnu_171_in_2, msg_to_bit_it_11_vnu_172_in_0, msg_to_bit_it_11_vnu_172_in_1, msg_to_bit_it_11_vnu_172_in_2, msg_to_bit_it_11_vnu_173_in_0, msg_to_bit_it_11_vnu_173_in_1, msg_to_bit_it_11_vnu_173_in_2, msg_to_bit_it_11_vnu_174_in_0, msg_to_bit_it_11_vnu_174_in_1, msg_to_bit_it_11_vnu_174_in_2, msg_to_bit_it_11_vnu_175_in_0, msg_to_bit_it_11_vnu_175_in_1, msg_to_bit_it_11_vnu_175_in_2, msg_to_bit_it_11_vnu_176_in_0, msg_to_bit_it_11_vnu_176_in_1, msg_to_bit_it_11_vnu_176_in_2, msg_to_bit_it_11_vnu_177_in_0, msg_to_bit_it_11_vnu_177_in_1, msg_to_bit_it_11_vnu_177_in_2, msg_to_bit_it_11_vnu_178_in_0, msg_to_bit_it_11_vnu_178_in_1, msg_to_bit_it_11_vnu_178_in_2, msg_to_bit_it_11_vnu_179_in_0, msg_to_bit_it_11_vnu_179_in_1, msg_to_bit_it_11_vnu_179_in_2, msg_to_bit_it_11_vnu_180_in_0, msg_to_bit_it_11_vnu_180_in_1, msg_to_bit_it_11_vnu_180_in_2, msg_to_bit_it_11_vnu_181_in_0, msg_to_bit_it_11_vnu_181_in_1, msg_to_bit_it_11_vnu_181_in_2, msg_to_bit_it_11_vnu_182_in_0, msg_to_bit_it_11_vnu_182_in_1, msg_to_bit_it_11_vnu_182_in_2, msg_to_bit_it_11_vnu_183_in_0, msg_to_bit_it_11_vnu_183_in_1, msg_to_bit_it_11_vnu_183_in_2, msg_to_bit_it_11_vnu_184_in_0, msg_to_bit_it_11_vnu_184_in_1, msg_to_bit_it_11_vnu_184_in_2, msg_to_bit_it_11_vnu_185_in_0, msg_to_bit_it_11_vnu_185_in_1, msg_to_bit_it_11_vnu_185_in_2, msg_to_bit_it_11_vnu_186_in_0, msg_to_bit_it_11_vnu_186_in_1, msg_to_bit_it_11_vnu_186_in_2, msg_to_bit_it_11_vnu_187_in_0, msg_to_bit_it_11_vnu_187_in_1, msg_to_bit_it_11_vnu_187_in_2, msg_to_bit_it_11_vnu_188_in_0, msg_to_bit_it_11_vnu_188_in_1, msg_to_bit_it_11_vnu_188_in_2, msg_to_bit_it_11_vnu_189_in_0, msg_to_bit_it_11_vnu_189_in_1, msg_to_bit_it_11_vnu_189_in_2, msg_to_bit_it_11_vnu_190_in_0, msg_to_bit_it_11_vnu_190_in_1, msg_to_bit_it_11_vnu_190_in_2, msg_to_bit_it_11_vnu_191_in_0, msg_to_bit_it_11_vnu_191_in_1, msg_to_bit_it_11_vnu_191_in_2, msg_to_bit_it_11_vnu_192_in_0, msg_to_bit_it_11_vnu_192_in_1, msg_to_bit_it_11_vnu_192_in_2, msg_to_bit_it_11_vnu_193_in_0, msg_to_bit_it_11_vnu_193_in_1, msg_to_bit_it_11_vnu_193_in_2, msg_to_bit_it_11_vnu_194_in_0, msg_to_bit_it_11_vnu_194_in_1, msg_to_bit_it_11_vnu_194_in_2, msg_to_bit_it_11_vnu_195_in_0, msg_to_bit_it_11_vnu_195_in_1, msg_to_bit_it_11_vnu_195_in_2, msg_to_bit_it_11_vnu_196_in_0, msg_to_bit_it_11_vnu_196_in_1, msg_to_bit_it_11_vnu_196_in_2, msg_to_bit_it_11_vnu_197_in_0, msg_to_bit_it_11_vnu_197_in_1, msg_to_bit_it_11_vnu_197_in_2, msg_to_bit_it_12_vnu_0_in_0, msg_to_bit_it_12_vnu_0_in_1, msg_to_bit_it_12_vnu_0_in_2, msg_to_bit_it_12_vnu_1_in_0, msg_to_bit_it_12_vnu_1_in_1, msg_to_bit_it_12_vnu_1_in_2, msg_to_bit_it_12_vnu_2_in_0, msg_to_bit_it_12_vnu_2_in_1, msg_to_bit_it_12_vnu_2_in_2, msg_to_bit_it_12_vnu_3_in_0, msg_to_bit_it_12_vnu_3_in_1, msg_to_bit_it_12_vnu_3_in_2, msg_to_bit_it_12_vnu_4_in_0, msg_to_bit_it_12_vnu_4_in_1, msg_to_bit_it_12_vnu_4_in_2, msg_to_bit_it_12_vnu_5_in_0, msg_to_bit_it_12_vnu_5_in_1, msg_to_bit_it_12_vnu_5_in_2, msg_to_bit_it_12_vnu_6_in_0, msg_to_bit_it_12_vnu_6_in_1, msg_to_bit_it_12_vnu_6_in_2, msg_to_bit_it_12_vnu_7_in_0, msg_to_bit_it_12_vnu_7_in_1, msg_to_bit_it_12_vnu_7_in_2, msg_to_bit_it_12_vnu_8_in_0, msg_to_bit_it_12_vnu_8_in_1, msg_to_bit_it_12_vnu_8_in_2, msg_to_bit_it_12_vnu_9_in_0, msg_to_bit_it_12_vnu_9_in_1, msg_to_bit_it_12_vnu_9_in_2, msg_to_bit_it_12_vnu_10_in_0, msg_to_bit_it_12_vnu_10_in_1, msg_to_bit_it_12_vnu_10_in_2, msg_to_bit_it_12_vnu_11_in_0, msg_to_bit_it_12_vnu_11_in_1, msg_to_bit_it_12_vnu_11_in_2, msg_to_bit_it_12_vnu_12_in_0, msg_to_bit_it_12_vnu_12_in_1, msg_to_bit_it_12_vnu_12_in_2, msg_to_bit_it_12_vnu_13_in_0, msg_to_bit_it_12_vnu_13_in_1, msg_to_bit_it_12_vnu_13_in_2, msg_to_bit_it_12_vnu_14_in_0, msg_to_bit_it_12_vnu_14_in_1, msg_to_bit_it_12_vnu_14_in_2, msg_to_bit_it_12_vnu_15_in_0, msg_to_bit_it_12_vnu_15_in_1, msg_to_bit_it_12_vnu_15_in_2, msg_to_bit_it_12_vnu_16_in_0, msg_to_bit_it_12_vnu_16_in_1, msg_to_bit_it_12_vnu_16_in_2, msg_to_bit_it_12_vnu_17_in_0, msg_to_bit_it_12_vnu_17_in_1, msg_to_bit_it_12_vnu_17_in_2, msg_to_bit_it_12_vnu_18_in_0, msg_to_bit_it_12_vnu_18_in_1, msg_to_bit_it_12_vnu_18_in_2, msg_to_bit_it_12_vnu_19_in_0, msg_to_bit_it_12_vnu_19_in_1, msg_to_bit_it_12_vnu_19_in_2, msg_to_bit_it_12_vnu_20_in_0, msg_to_bit_it_12_vnu_20_in_1, msg_to_bit_it_12_vnu_20_in_2, msg_to_bit_it_12_vnu_21_in_0, msg_to_bit_it_12_vnu_21_in_1, msg_to_bit_it_12_vnu_21_in_2, msg_to_bit_it_12_vnu_22_in_0, msg_to_bit_it_12_vnu_22_in_1, msg_to_bit_it_12_vnu_22_in_2, msg_to_bit_it_12_vnu_23_in_0, msg_to_bit_it_12_vnu_23_in_1, msg_to_bit_it_12_vnu_23_in_2, msg_to_bit_it_12_vnu_24_in_0, msg_to_bit_it_12_vnu_24_in_1, msg_to_bit_it_12_vnu_24_in_2, msg_to_bit_it_12_vnu_25_in_0, msg_to_bit_it_12_vnu_25_in_1, msg_to_bit_it_12_vnu_25_in_2, msg_to_bit_it_12_vnu_26_in_0, msg_to_bit_it_12_vnu_26_in_1, msg_to_bit_it_12_vnu_26_in_2, msg_to_bit_it_12_vnu_27_in_0, msg_to_bit_it_12_vnu_27_in_1, msg_to_bit_it_12_vnu_27_in_2, msg_to_bit_it_12_vnu_28_in_0, msg_to_bit_it_12_vnu_28_in_1, msg_to_bit_it_12_vnu_28_in_2, msg_to_bit_it_12_vnu_29_in_0, msg_to_bit_it_12_vnu_29_in_1, msg_to_bit_it_12_vnu_29_in_2, msg_to_bit_it_12_vnu_30_in_0, msg_to_bit_it_12_vnu_30_in_1, msg_to_bit_it_12_vnu_30_in_2, msg_to_bit_it_12_vnu_31_in_0, msg_to_bit_it_12_vnu_31_in_1, msg_to_bit_it_12_vnu_31_in_2, msg_to_bit_it_12_vnu_32_in_0, msg_to_bit_it_12_vnu_32_in_1, msg_to_bit_it_12_vnu_32_in_2, msg_to_bit_it_12_vnu_33_in_0, msg_to_bit_it_12_vnu_33_in_1, msg_to_bit_it_12_vnu_33_in_2, msg_to_bit_it_12_vnu_34_in_0, msg_to_bit_it_12_vnu_34_in_1, msg_to_bit_it_12_vnu_34_in_2, msg_to_bit_it_12_vnu_35_in_0, msg_to_bit_it_12_vnu_35_in_1, msg_to_bit_it_12_vnu_35_in_2, msg_to_bit_it_12_vnu_36_in_0, msg_to_bit_it_12_vnu_36_in_1, msg_to_bit_it_12_vnu_36_in_2, msg_to_bit_it_12_vnu_37_in_0, msg_to_bit_it_12_vnu_37_in_1, msg_to_bit_it_12_vnu_37_in_2, msg_to_bit_it_12_vnu_38_in_0, msg_to_bit_it_12_vnu_38_in_1, msg_to_bit_it_12_vnu_38_in_2, msg_to_bit_it_12_vnu_39_in_0, msg_to_bit_it_12_vnu_39_in_1, msg_to_bit_it_12_vnu_39_in_2, msg_to_bit_it_12_vnu_40_in_0, msg_to_bit_it_12_vnu_40_in_1, msg_to_bit_it_12_vnu_40_in_2, msg_to_bit_it_12_vnu_41_in_0, msg_to_bit_it_12_vnu_41_in_1, msg_to_bit_it_12_vnu_41_in_2, msg_to_bit_it_12_vnu_42_in_0, msg_to_bit_it_12_vnu_42_in_1, msg_to_bit_it_12_vnu_42_in_2, msg_to_bit_it_12_vnu_43_in_0, msg_to_bit_it_12_vnu_43_in_1, msg_to_bit_it_12_vnu_43_in_2, msg_to_bit_it_12_vnu_44_in_0, msg_to_bit_it_12_vnu_44_in_1, msg_to_bit_it_12_vnu_44_in_2, msg_to_bit_it_12_vnu_45_in_0, msg_to_bit_it_12_vnu_45_in_1, msg_to_bit_it_12_vnu_45_in_2, msg_to_bit_it_12_vnu_46_in_0, msg_to_bit_it_12_vnu_46_in_1, msg_to_bit_it_12_vnu_46_in_2, msg_to_bit_it_12_vnu_47_in_0, msg_to_bit_it_12_vnu_47_in_1, msg_to_bit_it_12_vnu_47_in_2, msg_to_bit_it_12_vnu_48_in_0, msg_to_bit_it_12_vnu_48_in_1, msg_to_bit_it_12_vnu_48_in_2, msg_to_bit_it_12_vnu_49_in_0, msg_to_bit_it_12_vnu_49_in_1, msg_to_bit_it_12_vnu_49_in_2, msg_to_bit_it_12_vnu_50_in_0, msg_to_bit_it_12_vnu_50_in_1, msg_to_bit_it_12_vnu_50_in_2, msg_to_bit_it_12_vnu_51_in_0, msg_to_bit_it_12_vnu_51_in_1, msg_to_bit_it_12_vnu_51_in_2, msg_to_bit_it_12_vnu_52_in_0, msg_to_bit_it_12_vnu_52_in_1, msg_to_bit_it_12_vnu_52_in_2, msg_to_bit_it_12_vnu_53_in_0, msg_to_bit_it_12_vnu_53_in_1, msg_to_bit_it_12_vnu_53_in_2, msg_to_bit_it_12_vnu_54_in_0, msg_to_bit_it_12_vnu_54_in_1, msg_to_bit_it_12_vnu_54_in_2, msg_to_bit_it_12_vnu_55_in_0, msg_to_bit_it_12_vnu_55_in_1, msg_to_bit_it_12_vnu_55_in_2, msg_to_bit_it_12_vnu_56_in_0, msg_to_bit_it_12_vnu_56_in_1, msg_to_bit_it_12_vnu_56_in_2, msg_to_bit_it_12_vnu_57_in_0, msg_to_bit_it_12_vnu_57_in_1, msg_to_bit_it_12_vnu_57_in_2, msg_to_bit_it_12_vnu_58_in_0, msg_to_bit_it_12_vnu_58_in_1, msg_to_bit_it_12_vnu_58_in_2, msg_to_bit_it_12_vnu_59_in_0, msg_to_bit_it_12_vnu_59_in_1, msg_to_bit_it_12_vnu_59_in_2, msg_to_bit_it_12_vnu_60_in_0, msg_to_bit_it_12_vnu_60_in_1, msg_to_bit_it_12_vnu_60_in_2, msg_to_bit_it_12_vnu_61_in_0, msg_to_bit_it_12_vnu_61_in_1, msg_to_bit_it_12_vnu_61_in_2, msg_to_bit_it_12_vnu_62_in_0, msg_to_bit_it_12_vnu_62_in_1, msg_to_bit_it_12_vnu_62_in_2, msg_to_bit_it_12_vnu_63_in_0, msg_to_bit_it_12_vnu_63_in_1, msg_to_bit_it_12_vnu_63_in_2, msg_to_bit_it_12_vnu_64_in_0, msg_to_bit_it_12_vnu_64_in_1, msg_to_bit_it_12_vnu_64_in_2, msg_to_bit_it_12_vnu_65_in_0, msg_to_bit_it_12_vnu_65_in_1, msg_to_bit_it_12_vnu_65_in_2, msg_to_bit_it_12_vnu_66_in_0, msg_to_bit_it_12_vnu_66_in_1, msg_to_bit_it_12_vnu_66_in_2, msg_to_bit_it_12_vnu_67_in_0, msg_to_bit_it_12_vnu_67_in_1, msg_to_bit_it_12_vnu_67_in_2, msg_to_bit_it_12_vnu_68_in_0, msg_to_bit_it_12_vnu_68_in_1, msg_to_bit_it_12_vnu_68_in_2, msg_to_bit_it_12_vnu_69_in_0, msg_to_bit_it_12_vnu_69_in_1, msg_to_bit_it_12_vnu_69_in_2, msg_to_bit_it_12_vnu_70_in_0, msg_to_bit_it_12_vnu_70_in_1, msg_to_bit_it_12_vnu_70_in_2, msg_to_bit_it_12_vnu_71_in_0, msg_to_bit_it_12_vnu_71_in_1, msg_to_bit_it_12_vnu_71_in_2, msg_to_bit_it_12_vnu_72_in_0, msg_to_bit_it_12_vnu_72_in_1, msg_to_bit_it_12_vnu_72_in_2, msg_to_bit_it_12_vnu_73_in_0, msg_to_bit_it_12_vnu_73_in_1, msg_to_bit_it_12_vnu_73_in_2, msg_to_bit_it_12_vnu_74_in_0, msg_to_bit_it_12_vnu_74_in_1, msg_to_bit_it_12_vnu_74_in_2, msg_to_bit_it_12_vnu_75_in_0, msg_to_bit_it_12_vnu_75_in_1, msg_to_bit_it_12_vnu_75_in_2, msg_to_bit_it_12_vnu_76_in_0, msg_to_bit_it_12_vnu_76_in_1, msg_to_bit_it_12_vnu_76_in_2, msg_to_bit_it_12_vnu_77_in_0, msg_to_bit_it_12_vnu_77_in_1, msg_to_bit_it_12_vnu_77_in_2, msg_to_bit_it_12_vnu_78_in_0, msg_to_bit_it_12_vnu_78_in_1, msg_to_bit_it_12_vnu_78_in_2, msg_to_bit_it_12_vnu_79_in_0, msg_to_bit_it_12_vnu_79_in_1, msg_to_bit_it_12_vnu_79_in_2, msg_to_bit_it_12_vnu_80_in_0, msg_to_bit_it_12_vnu_80_in_1, msg_to_bit_it_12_vnu_80_in_2, msg_to_bit_it_12_vnu_81_in_0, msg_to_bit_it_12_vnu_81_in_1, msg_to_bit_it_12_vnu_81_in_2, msg_to_bit_it_12_vnu_82_in_0, msg_to_bit_it_12_vnu_82_in_1, msg_to_bit_it_12_vnu_82_in_2, msg_to_bit_it_12_vnu_83_in_0, msg_to_bit_it_12_vnu_83_in_1, msg_to_bit_it_12_vnu_83_in_2, msg_to_bit_it_12_vnu_84_in_0, msg_to_bit_it_12_vnu_84_in_1, msg_to_bit_it_12_vnu_84_in_2, msg_to_bit_it_12_vnu_85_in_0, msg_to_bit_it_12_vnu_85_in_1, msg_to_bit_it_12_vnu_85_in_2, msg_to_bit_it_12_vnu_86_in_0, msg_to_bit_it_12_vnu_86_in_1, msg_to_bit_it_12_vnu_86_in_2, msg_to_bit_it_12_vnu_87_in_0, msg_to_bit_it_12_vnu_87_in_1, msg_to_bit_it_12_vnu_87_in_2, msg_to_bit_it_12_vnu_88_in_0, msg_to_bit_it_12_vnu_88_in_1, msg_to_bit_it_12_vnu_88_in_2, msg_to_bit_it_12_vnu_89_in_0, msg_to_bit_it_12_vnu_89_in_1, msg_to_bit_it_12_vnu_89_in_2, msg_to_bit_it_12_vnu_90_in_0, msg_to_bit_it_12_vnu_90_in_1, msg_to_bit_it_12_vnu_90_in_2, msg_to_bit_it_12_vnu_91_in_0, msg_to_bit_it_12_vnu_91_in_1, msg_to_bit_it_12_vnu_91_in_2, msg_to_bit_it_12_vnu_92_in_0, msg_to_bit_it_12_vnu_92_in_1, msg_to_bit_it_12_vnu_92_in_2, msg_to_bit_it_12_vnu_93_in_0, msg_to_bit_it_12_vnu_93_in_1, msg_to_bit_it_12_vnu_93_in_2, msg_to_bit_it_12_vnu_94_in_0, msg_to_bit_it_12_vnu_94_in_1, msg_to_bit_it_12_vnu_94_in_2, msg_to_bit_it_12_vnu_95_in_0, msg_to_bit_it_12_vnu_95_in_1, msg_to_bit_it_12_vnu_95_in_2, msg_to_bit_it_12_vnu_96_in_0, msg_to_bit_it_12_vnu_96_in_1, msg_to_bit_it_12_vnu_96_in_2, msg_to_bit_it_12_vnu_97_in_0, msg_to_bit_it_12_vnu_97_in_1, msg_to_bit_it_12_vnu_97_in_2, msg_to_bit_it_12_vnu_98_in_0, msg_to_bit_it_12_vnu_98_in_1, msg_to_bit_it_12_vnu_98_in_2, msg_to_bit_it_12_vnu_99_in_0, msg_to_bit_it_12_vnu_99_in_1, msg_to_bit_it_12_vnu_99_in_2, msg_to_bit_it_12_vnu_100_in_0, msg_to_bit_it_12_vnu_100_in_1, msg_to_bit_it_12_vnu_100_in_2, msg_to_bit_it_12_vnu_101_in_0, msg_to_bit_it_12_vnu_101_in_1, msg_to_bit_it_12_vnu_101_in_2, msg_to_bit_it_12_vnu_102_in_0, msg_to_bit_it_12_vnu_102_in_1, msg_to_bit_it_12_vnu_102_in_2, msg_to_bit_it_12_vnu_103_in_0, msg_to_bit_it_12_vnu_103_in_1, msg_to_bit_it_12_vnu_103_in_2, msg_to_bit_it_12_vnu_104_in_0, msg_to_bit_it_12_vnu_104_in_1, msg_to_bit_it_12_vnu_104_in_2, msg_to_bit_it_12_vnu_105_in_0, msg_to_bit_it_12_vnu_105_in_1, msg_to_bit_it_12_vnu_105_in_2, msg_to_bit_it_12_vnu_106_in_0, msg_to_bit_it_12_vnu_106_in_1, msg_to_bit_it_12_vnu_106_in_2, msg_to_bit_it_12_vnu_107_in_0, msg_to_bit_it_12_vnu_107_in_1, msg_to_bit_it_12_vnu_107_in_2, msg_to_bit_it_12_vnu_108_in_0, msg_to_bit_it_12_vnu_108_in_1, msg_to_bit_it_12_vnu_108_in_2, msg_to_bit_it_12_vnu_109_in_0, msg_to_bit_it_12_vnu_109_in_1, msg_to_bit_it_12_vnu_109_in_2, msg_to_bit_it_12_vnu_110_in_0, msg_to_bit_it_12_vnu_110_in_1, msg_to_bit_it_12_vnu_110_in_2, msg_to_bit_it_12_vnu_111_in_0, msg_to_bit_it_12_vnu_111_in_1, msg_to_bit_it_12_vnu_111_in_2, msg_to_bit_it_12_vnu_112_in_0, msg_to_bit_it_12_vnu_112_in_1, msg_to_bit_it_12_vnu_112_in_2, msg_to_bit_it_12_vnu_113_in_0, msg_to_bit_it_12_vnu_113_in_1, msg_to_bit_it_12_vnu_113_in_2, msg_to_bit_it_12_vnu_114_in_0, msg_to_bit_it_12_vnu_114_in_1, msg_to_bit_it_12_vnu_114_in_2, msg_to_bit_it_12_vnu_115_in_0, msg_to_bit_it_12_vnu_115_in_1, msg_to_bit_it_12_vnu_115_in_2, msg_to_bit_it_12_vnu_116_in_0, msg_to_bit_it_12_vnu_116_in_1, msg_to_bit_it_12_vnu_116_in_2, msg_to_bit_it_12_vnu_117_in_0, msg_to_bit_it_12_vnu_117_in_1, msg_to_bit_it_12_vnu_117_in_2, msg_to_bit_it_12_vnu_118_in_0, msg_to_bit_it_12_vnu_118_in_1, msg_to_bit_it_12_vnu_118_in_2, msg_to_bit_it_12_vnu_119_in_0, msg_to_bit_it_12_vnu_119_in_1, msg_to_bit_it_12_vnu_119_in_2, msg_to_bit_it_12_vnu_120_in_0, msg_to_bit_it_12_vnu_120_in_1, msg_to_bit_it_12_vnu_120_in_2, msg_to_bit_it_12_vnu_121_in_0, msg_to_bit_it_12_vnu_121_in_1, msg_to_bit_it_12_vnu_121_in_2, msg_to_bit_it_12_vnu_122_in_0, msg_to_bit_it_12_vnu_122_in_1, msg_to_bit_it_12_vnu_122_in_2, msg_to_bit_it_12_vnu_123_in_0, msg_to_bit_it_12_vnu_123_in_1, msg_to_bit_it_12_vnu_123_in_2, msg_to_bit_it_12_vnu_124_in_0, msg_to_bit_it_12_vnu_124_in_1, msg_to_bit_it_12_vnu_124_in_2, msg_to_bit_it_12_vnu_125_in_0, msg_to_bit_it_12_vnu_125_in_1, msg_to_bit_it_12_vnu_125_in_2, msg_to_bit_it_12_vnu_126_in_0, msg_to_bit_it_12_vnu_126_in_1, msg_to_bit_it_12_vnu_126_in_2, msg_to_bit_it_12_vnu_127_in_0, msg_to_bit_it_12_vnu_127_in_1, msg_to_bit_it_12_vnu_127_in_2, msg_to_bit_it_12_vnu_128_in_0, msg_to_bit_it_12_vnu_128_in_1, msg_to_bit_it_12_vnu_128_in_2, msg_to_bit_it_12_vnu_129_in_0, msg_to_bit_it_12_vnu_129_in_1, msg_to_bit_it_12_vnu_129_in_2, msg_to_bit_it_12_vnu_130_in_0, msg_to_bit_it_12_vnu_130_in_1, msg_to_bit_it_12_vnu_130_in_2, msg_to_bit_it_12_vnu_131_in_0, msg_to_bit_it_12_vnu_131_in_1, msg_to_bit_it_12_vnu_131_in_2, msg_to_bit_it_12_vnu_132_in_0, msg_to_bit_it_12_vnu_132_in_1, msg_to_bit_it_12_vnu_132_in_2, msg_to_bit_it_12_vnu_133_in_0, msg_to_bit_it_12_vnu_133_in_1, msg_to_bit_it_12_vnu_133_in_2, msg_to_bit_it_12_vnu_134_in_0, msg_to_bit_it_12_vnu_134_in_1, msg_to_bit_it_12_vnu_134_in_2, msg_to_bit_it_12_vnu_135_in_0, msg_to_bit_it_12_vnu_135_in_1, msg_to_bit_it_12_vnu_135_in_2, msg_to_bit_it_12_vnu_136_in_0, msg_to_bit_it_12_vnu_136_in_1, msg_to_bit_it_12_vnu_136_in_2, msg_to_bit_it_12_vnu_137_in_0, msg_to_bit_it_12_vnu_137_in_1, msg_to_bit_it_12_vnu_137_in_2, msg_to_bit_it_12_vnu_138_in_0, msg_to_bit_it_12_vnu_138_in_1, msg_to_bit_it_12_vnu_138_in_2, msg_to_bit_it_12_vnu_139_in_0, msg_to_bit_it_12_vnu_139_in_1, msg_to_bit_it_12_vnu_139_in_2, msg_to_bit_it_12_vnu_140_in_0, msg_to_bit_it_12_vnu_140_in_1, msg_to_bit_it_12_vnu_140_in_2, msg_to_bit_it_12_vnu_141_in_0, msg_to_bit_it_12_vnu_141_in_1, msg_to_bit_it_12_vnu_141_in_2, msg_to_bit_it_12_vnu_142_in_0, msg_to_bit_it_12_vnu_142_in_1, msg_to_bit_it_12_vnu_142_in_2, msg_to_bit_it_12_vnu_143_in_0, msg_to_bit_it_12_vnu_143_in_1, msg_to_bit_it_12_vnu_143_in_2, msg_to_bit_it_12_vnu_144_in_0, msg_to_bit_it_12_vnu_144_in_1, msg_to_bit_it_12_vnu_144_in_2, msg_to_bit_it_12_vnu_145_in_0, msg_to_bit_it_12_vnu_145_in_1, msg_to_bit_it_12_vnu_145_in_2, msg_to_bit_it_12_vnu_146_in_0, msg_to_bit_it_12_vnu_146_in_1, msg_to_bit_it_12_vnu_146_in_2, msg_to_bit_it_12_vnu_147_in_0, msg_to_bit_it_12_vnu_147_in_1, msg_to_bit_it_12_vnu_147_in_2, msg_to_bit_it_12_vnu_148_in_0, msg_to_bit_it_12_vnu_148_in_1, msg_to_bit_it_12_vnu_148_in_2, msg_to_bit_it_12_vnu_149_in_0, msg_to_bit_it_12_vnu_149_in_1, msg_to_bit_it_12_vnu_149_in_2, msg_to_bit_it_12_vnu_150_in_0, msg_to_bit_it_12_vnu_150_in_1, msg_to_bit_it_12_vnu_150_in_2, msg_to_bit_it_12_vnu_151_in_0, msg_to_bit_it_12_vnu_151_in_1, msg_to_bit_it_12_vnu_151_in_2, msg_to_bit_it_12_vnu_152_in_0, msg_to_bit_it_12_vnu_152_in_1, msg_to_bit_it_12_vnu_152_in_2, msg_to_bit_it_12_vnu_153_in_0, msg_to_bit_it_12_vnu_153_in_1, msg_to_bit_it_12_vnu_153_in_2, msg_to_bit_it_12_vnu_154_in_0, msg_to_bit_it_12_vnu_154_in_1, msg_to_bit_it_12_vnu_154_in_2, msg_to_bit_it_12_vnu_155_in_0, msg_to_bit_it_12_vnu_155_in_1, msg_to_bit_it_12_vnu_155_in_2, msg_to_bit_it_12_vnu_156_in_0, msg_to_bit_it_12_vnu_156_in_1, msg_to_bit_it_12_vnu_156_in_2, msg_to_bit_it_12_vnu_157_in_0, msg_to_bit_it_12_vnu_157_in_1, msg_to_bit_it_12_vnu_157_in_2, msg_to_bit_it_12_vnu_158_in_0, msg_to_bit_it_12_vnu_158_in_1, msg_to_bit_it_12_vnu_158_in_2, msg_to_bit_it_12_vnu_159_in_0, msg_to_bit_it_12_vnu_159_in_1, msg_to_bit_it_12_vnu_159_in_2, msg_to_bit_it_12_vnu_160_in_0, msg_to_bit_it_12_vnu_160_in_1, msg_to_bit_it_12_vnu_160_in_2, msg_to_bit_it_12_vnu_161_in_0, msg_to_bit_it_12_vnu_161_in_1, msg_to_bit_it_12_vnu_161_in_2, msg_to_bit_it_12_vnu_162_in_0, msg_to_bit_it_12_vnu_162_in_1, msg_to_bit_it_12_vnu_162_in_2, msg_to_bit_it_12_vnu_163_in_0, msg_to_bit_it_12_vnu_163_in_1, msg_to_bit_it_12_vnu_163_in_2, msg_to_bit_it_12_vnu_164_in_0, msg_to_bit_it_12_vnu_164_in_1, msg_to_bit_it_12_vnu_164_in_2, msg_to_bit_it_12_vnu_165_in_0, msg_to_bit_it_12_vnu_165_in_1, msg_to_bit_it_12_vnu_165_in_2, msg_to_bit_it_12_vnu_166_in_0, msg_to_bit_it_12_vnu_166_in_1, msg_to_bit_it_12_vnu_166_in_2, msg_to_bit_it_12_vnu_167_in_0, msg_to_bit_it_12_vnu_167_in_1, msg_to_bit_it_12_vnu_167_in_2, msg_to_bit_it_12_vnu_168_in_0, msg_to_bit_it_12_vnu_168_in_1, msg_to_bit_it_12_vnu_168_in_2, msg_to_bit_it_12_vnu_169_in_0, msg_to_bit_it_12_vnu_169_in_1, msg_to_bit_it_12_vnu_169_in_2, msg_to_bit_it_12_vnu_170_in_0, msg_to_bit_it_12_vnu_170_in_1, msg_to_bit_it_12_vnu_170_in_2, msg_to_bit_it_12_vnu_171_in_0, msg_to_bit_it_12_vnu_171_in_1, msg_to_bit_it_12_vnu_171_in_2, msg_to_bit_it_12_vnu_172_in_0, msg_to_bit_it_12_vnu_172_in_1, msg_to_bit_it_12_vnu_172_in_2, msg_to_bit_it_12_vnu_173_in_0, msg_to_bit_it_12_vnu_173_in_1, msg_to_bit_it_12_vnu_173_in_2, msg_to_bit_it_12_vnu_174_in_0, msg_to_bit_it_12_vnu_174_in_1, msg_to_bit_it_12_vnu_174_in_2, msg_to_bit_it_12_vnu_175_in_0, msg_to_bit_it_12_vnu_175_in_1, msg_to_bit_it_12_vnu_175_in_2, msg_to_bit_it_12_vnu_176_in_0, msg_to_bit_it_12_vnu_176_in_1, msg_to_bit_it_12_vnu_176_in_2, msg_to_bit_it_12_vnu_177_in_0, msg_to_bit_it_12_vnu_177_in_1, msg_to_bit_it_12_vnu_177_in_2, msg_to_bit_it_12_vnu_178_in_0, msg_to_bit_it_12_vnu_178_in_1, msg_to_bit_it_12_vnu_178_in_2, msg_to_bit_it_12_vnu_179_in_0, msg_to_bit_it_12_vnu_179_in_1, msg_to_bit_it_12_vnu_179_in_2, msg_to_bit_it_12_vnu_180_in_0, msg_to_bit_it_12_vnu_180_in_1, msg_to_bit_it_12_vnu_180_in_2, msg_to_bit_it_12_vnu_181_in_0, msg_to_bit_it_12_vnu_181_in_1, msg_to_bit_it_12_vnu_181_in_2, msg_to_bit_it_12_vnu_182_in_0, msg_to_bit_it_12_vnu_182_in_1, msg_to_bit_it_12_vnu_182_in_2, msg_to_bit_it_12_vnu_183_in_0, msg_to_bit_it_12_vnu_183_in_1, msg_to_bit_it_12_vnu_183_in_2, msg_to_bit_it_12_vnu_184_in_0, msg_to_bit_it_12_vnu_184_in_1, msg_to_bit_it_12_vnu_184_in_2, msg_to_bit_it_12_vnu_185_in_0, msg_to_bit_it_12_vnu_185_in_1, msg_to_bit_it_12_vnu_185_in_2, msg_to_bit_it_12_vnu_186_in_0, msg_to_bit_it_12_vnu_186_in_1, msg_to_bit_it_12_vnu_186_in_2, msg_to_bit_it_12_vnu_187_in_0, msg_to_bit_it_12_vnu_187_in_1, msg_to_bit_it_12_vnu_187_in_2, msg_to_bit_it_12_vnu_188_in_0, msg_to_bit_it_12_vnu_188_in_1, msg_to_bit_it_12_vnu_188_in_2, msg_to_bit_it_12_vnu_189_in_0, msg_to_bit_it_12_vnu_189_in_1, msg_to_bit_it_12_vnu_189_in_2, msg_to_bit_it_12_vnu_190_in_0, msg_to_bit_it_12_vnu_190_in_1, msg_to_bit_it_12_vnu_190_in_2, msg_to_bit_it_12_vnu_191_in_0, msg_to_bit_it_12_vnu_191_in_1, msg_to_bit_it_12_vnu_191_in_2, msg_to_bit_it_12_vnu_192_in_0, msg_to_bit_it_12_vnu_192_in_1, msg_to_bit_it_12_vnu_192_in_2, msg_to_bit_it_12_vnu_193_in_0, msg_to_bit_it_12_vnu_193_in_1, msg_to_bit_it_12_vnu_193_in_2, msg_to_bit_it_12_vnu_194_in_0, msg_to_bit_it_12_vnu_194_in_1, msg_to_bit_it_12_vnu_194_in_2, msg_to_bit_it_12_vnu_195_in_0, msg_to_bit_it_12_vnu_195_in_1, msg_to_bit_it_12_vnu_195_in_2, msg_to_bit_it_12_vnu_196_in_0, msg_to_bit_it_12_vnu_196_in_1, msg_to_bit_it_12_vnu_196_in_2, msg_to_bit_it_12_vnu_197_in_0, msg_to_bit_it_12_vnu_197_in_1, msg_to_bit_it_12_vnu_197_in_2, msg_to_bit_it_13_vnu_0_in_0, msg_to_bit_it_13_vnu_0_in_1, msg_to_bit_it_13_vnu_0_in_2, msg_to_bit_it_13_vnu_1_in_0, msg_to_bit_it_13_vnu_1_in_1, msg_to_bit_it_13_vnu_1_in_2, msg_to_bit_it_13_vnu_2_in_0, msg_to_bit_it_13_vnu_2_in_1, msg_to_bit_it_13_vnu_2_in_2, msg_to_bit_it_13_vnu_3_in_0, msg_to_bit_it_13_vnu_3_in_1, msg_to_bit_it_13_vnu_3_in_2, msg_to_bit_it_13_vnu_4_in_0, msg_to_bit_it_13_vnu_4_in_1, msg_to_bit_it_13_vnu_4_in_2, msg_to_bit_it_13_vnu_5_in_0, msg_to_bit_it_13_vnu_5_in_1, msg_to_bit_it_13_vnu_5_in_2, msg_to_bit_it_13_vnu_6_in_0, msg_to_bit_it_13_vnu_6_in_1, msg_to_bit_it_13_vnu_6_in_2, msg_to_bit_it_13_vnu_7_in_0, msg_to_bit_it_13_vnu_7_in_1, msg_to_bit_it_13_vnu_7_in_2, msg_to_bit_it_13_vnu_8_in_0, msg_to_bit_it_13_vnu_8_in_1, msg_to_bit_it_13_vnu_8_in_2, msg_to_bit_it_13_vnu_9_in_0, msg_to_bit_it_13_vnu_9_in_1, msg_to_bit_it_13_vnu_9_in_2, msg_to_bit_it_13_vnu_10_in_0, msg_to_bit_it_13_vnu_10_in_1, msg_to_bit_it_13_vnu_10_in_2, msg_to_bit_it_13_vnu_11_in_0, msg_to_bit_it_13_vnu_11_in_1, msg_to_bit_it_13_vnu_11_in_2, msg_to_bit_it_13_vnu_12_in_0, msg_to_bit_it_13_vnu_12_in_1, msg_to_bit_it_13_vnu_12_in_2, msg_to_bit_it_13_vnu_13_in_0, msg_to_bit_it_13_vnu_13_in_1, msg_to_bit_it_13_vnu_13_in_2, msg_to_bit_it_13_vnu_14_in_0, msg_to_bit_it_13_vnu_14_in_1, msg_to_bit_it_13_vnu_14_in_2, msg_to_bit_it_13_vnu_15_in_0, msg_to_bit_it_13_vnu_15_in_1, msg_to_bit_it_13_vnu_15_in_2, msg_to_bit_it_13_vnu_16_in_0, msg_to_bit_it_13_vnu_16_in_1, msg_to_bit_it_13_vnu_16_in_2, msg_to_bit_it_13_vnu_17_in_0, msg_to_bit_it_13_vnu_17_in_1, msg_to_bit_it_13_vnu_17_in_2, msg_to_bit_it_13_vnu_18_in_0, msg_to_bit_it_13_vnu_18_in_1, msg_to_bit_it_13_vnu_18_in_2, msg_to_bit_it_13_vnu_19_in_0, msg_to_bit_it_13_vnu_19_in_1, msg_to_bit_it_13_vnu_19_in_2, msg_to_bit_it_13_vnu_20_in_0, msg_to_bit_it_13_vnu_20_in_1, msg_to_bit_it_13_vnu_20_in_2, msg_to_bit_it_13_vnu_21_in_0, msg_to_bit_it_13_vnu_21_in_1, msg_to_bit_it_13_vnu_21_in_2, msg_to_bit_it_13_vnu_22_in_0, msg_to_bit_it_13_vnu_22_in_1, msg_to_bit_it_13_vnu_22_in_2, msg_to_bit_it_13_vnu_23_in_0, msg_to_bit_it_13_vnu_23_in_1, msg_to_bit_it_13_vnu_23_in_2, msg_to_bit_it_13_vnu_24_in_0, msg_to_bit_it_13_vnu_24_in_1, msg_to_bit_it_13_vnu_24_in_2, msg_to_bit_it_13_vnu_25_in_0, msg_to_bit_it_13_vnu_25_in_1, msg_to_bit_it_13_vnu_25_in_2, msg_to_bit_it_13_vnu_26_in_0, msg_to_bit_it_13_vnu_26_in_1, msg_to_bit_it_13_vnu_26_in_2, msg_to_bit_it_13_vnu_27_in_0, msg_to_bit_it_13_vnu_27_in_1, msg_to_bit_it_13_vnu_27_in_2, msg_to_bit_it_13_vnu_28_in_0, msg_to_bit_it_13_vnu_28_in_1, msg_to_bit_it_13_vnu_28_in_2, msg_to_bit_it_13_vnu_29_in_0, msg_to_bit_it_13_vnu_29_in_1, msg_to_bit_it_13_vnu_29_in_2, msg_to_bit_it_13_vnu_30_in_0, msg_to_bit_it_13_vnu_30_in_1, msg_to_bit_it_13_vnu_30_in_2, msg_to_bit_it_13_vnu_31_in_0, msg_to_bit_it_13_vnu_31_in_1, msg_to_bit_it_13_vnu_31_in_2, msg_to_bit_it_13_vnu_32_in_0, msg_to_bit_it_13_vnu_32_in_1, msg_to_bit_it_13_vnu_32_in_2, msg_to_bit_it_13_vnu_33_in_0, msg_to_bit_it_13_vnu_33_in_1, msg_to_bit_it_13_vnu_33_in_2, msg_to_bit_it_13_vnu_34_in_0, msg_to_bit_it_13_vnu_34_in_1, msg_to_bit_it_13_vnu_34_in_2, msg_to_bit_it_13_vnu_35_in_0, msg_to_bit_it_13_vnu_35_in_1, msg_to_bit_it_13_vnu_35_in_2, msg_to_bit_it_13_vnu_36_in_0, msg_to_bit_it_13_vnu_36_in_1, msg_to_bit_it_13_vnu_36_in_2, msg_to_bit_it_13_vnu_37_in_0, msg_to_bit_it_13_vnu_37_in_1, msg_to_bit_it_13_vnu_37_in_2, msg_to_bit_it_13_vnu_38_in_0, msg_to_bit_it_13_vnu_38_in_1, msg_to_bit_it_13_vnu_38_in_2, msg_to_bit_it_13_vnu_39_in_0, msg_to_bit_it_13_vnu_39_in_1, msg_to_bit_it_13_vnu_39_in_2, msg_to_bit_it_13_vnu_40_in_0, msg_to_bit_it_13_vnu_40_in_1, msg_to_bit_it_13_vnu_40_in_2, msg_to_bit_it_13_vnu_41_in_0, msg_to_bit_it_13_vnu_41_in_1, msg_to_bit_it_13_vnu_41_in_2, msg_to_bit_it_13_vnu_42_in_0, msg_to_bit_it_13_vnu_42_in_1, msg_to_bit_it_13_vnu_42_in_2, msg_to_bit_it_13_vnu_43_in_0, msg_to_bit_it_13_vnu_43_in_1, msg_to_bit_it_13_vnu_43_in_2, msg_to_bit_it_13_vnu_44_in_0, msg_to_bit_it_13_vnu_44_in_1, msg_to_bit_it_13_vnu_44_in_2, msg_to_bit_it_13_vnu_45_in_0, msg_to_bit_it_13_vnu_45_in_1, msg_to_bit_it_13_vnu_45_in_2, msg_to_bit_it_13_vnu_46_in_0, msg_to_bit_it_13_vnu_46_in_1, msg_to_bit_it_13_vnu_46_in_2, msg_to_bit_it_13_vnu_47_in_0, msg_to_bit_it_13_vnu_47_in_1, msg_to_bit_it_13_vnu_47_in_2, msg_to_bit_it_13_vnu_48_in_0, msg_to_bit_it_13_vnu_48_in_1, msg_to_bit_it_13_vnu_48_in_2, msg_to_bit_it_13_vnu_49_in_0, msg_to_bit_it_13_vnu_49_in_1, msg_to_bit_it_13_vnu_49_in_2, msg_to_bit_it_13_vnu_50_in_0, msg_to_bit_it_13_vnu_50_in_1, msg_to_bit_it_13_vnu_50_in_2, msg_to_bit_it_13_vnu_51_in_0, msg_to_bit_it_13_vnu_51_in_1, msg_to_bit_it_13_vnu_51_in_2, msg_to_bit_it_13_vnu_52_in_0, msg_to_bit_it_13_vnu_52_in_1, msg_to_bit_it_13_vnu_52_in_2, msg_to_bit_it_13_vnu_53_in_0, msg_to_bit_it_13_vnu_53_in_1, msg_to_bit_it_13_vnu_53_in_2, msg_to_bit_it_13_vnu_54_in_0, msg_to_bit_it_13_vnu_54_in_1, msg_to_bit_it_13_vnu_54_in_2, msg_to_bit_it_13_vnu_55_in_0, msg_to_bit_it_13_vnu_55_in_1, msg_to_bit_it_13_vnu_55_in_2, msg_to_bit_it_13_vnu_56_in_0, msg_to_bit_it_13_vnu_56_in_1, msg_to_bit_it_13_vnu_56_in_2, msg_to_bit_it_13_vnu_57_in_0, msg_to_bit_it_13_vnu_57_in_1, msg_to_bit_it_13_vnu_57_in_2, msg_to_bit_it_13_vnu_58_in_0, msg_to_bit_it_13_vnu_58_in_1, msg_to_bit_it_13_vnu_58_in_2, msg_to_bit_it_13_vnu_59_in_0, msg_to_bit_it_13_vnu_59_in_1, msg_to_bit_it_13_vnu_59_in_2, msg_to_bit_it_13_vnu_60_in_0, msg_to_bit_it_13_vnu_60_in_1, msg_to_bit_it_13_vnu_60_in_2, msg_to_bit_it_13_vnu_61_in_0, msg_to_bit_it_13_vnu_61_in_1, msg_to_bit_it_13_vnu_61_in_2, msg_to_bit_it_13_vnu_62_in_0, msg_to_bit_it_13_vnu_62_in_1, msg_to_bit_it_13_vnu_62_in_2, msg_to_bit_it_13_vnu_63_in_0, msg_to_bit_it_13_vnu_63_in_1, msg_to_bit_it_13_vnu_63_in_2, msg_to_bit_it_13_vnu_64_in_0, msg_to_bit_it_13_vnu_64_in_1, msg_to_bit_it_13_vnu_64_in_2, msg_to_bit_it_13_vnu_65_in_0, msg_to_bit_it_13_vnu_65_in_1, msg_to_bit_it_13_vnu_65_in_2, msg_to_bit_it_13_vnu_66_in_0, msg_to_bit_it_13_vnu_66_in_1, msg_to_bit_it_13_vnu_66_in_2, msg_to_bit_it_13_vnu_67_in_0, msg_to_bit_it_13_vnu_67_in_1, msg_to_bit_it_13_vnu_67_in_2, msg_to_bit_it_13_vnu_68_in_0, msg_to_bit_it_13_vnu_68_in_1, msg_to_bit_it_13_vnu_68_in_2, msg_to_bit_it_13_vnu_69_in_0, msg_to_bit_it_13_vnu_69_in_1, msg_to_bit_it_13_vnu_69_in_2, msg_to_bit_it_13_vnu_70_in_0, msg_to_bit_it_13_vnu_70_in_1, msg_to_bit_it_13_vnu_70_in_2, msg_to_bit_it_13_vnu_71_in_0, msg_to_bit_it_13_vnu_71_in_1, msg_to_bit_it_13_vnu_71_in_2, msg_to_bit_it_13_vnu_72_in_0, msg_to_bit_it_13_vnu_72_in_1, msg_to_bit_it_13_vnu_72_in_2, msg_to_bit_it_13_vnu_73_in_0, msg_to_bit_it_13_vnu_73_in_1, msg_to_bit_it_13_vnu_73_in_2, msg_to_bit_it_13_vnu_74_in_0, msg_to_bit_it_13_vnu_74_in_1, msg_to_bit_it_13_vnu_74_in_2, msg_to_bit_it_13_vnu_75_in_0, msg_to_bit_it_13_vnu_75_in_1, msg_to_bit_it_13_vnu_75_in_2, msg_to_bit_it_13_vnu_76_in_0, msg_to_bit_it_13_vnu_76_in_1, msg_to_bit_it_13_vnu_76_in_2, msg_to_bit_it_13_vnu_77_in_0, msg_to_bit_it_13_vnu_77_in_1, msg_to_bit_it_13_vnu_77_in_2, msg_to_bit_it_13_vnu_78_in_0, msg_to_bit_it_13_vnu_78_in_1, msg_to_bit_it_13_vnu_78_in_2, msg_to_bit_it_13_vnu_79_in_0, msg_to_bit_it_13_vnu_79_in_1, msg_to_bit_it_13_vnu_79_in_2, msg_to_bit_it_13_vnu_80_in_0, msg_to_bit_it_13_vnu_80_in_1, msg_to_bit_it_13_vnu_80_in_2, msg_to_bit_it_13_vnu_81_in_0, msg_to_bit_it_13_vnu_81_in_1, msg_to_bit_it_13_vnu_81_in_2, msg_to_bit_it_13_vnu_82_in_0, msg_to_bit_it_13_vnu_82_in_1, msg_to_bit_it_13_vnu_82_in_2, msg_to_bit_it_13_vnu_83_in_0, msg_to_bit_it_13_vnu_83_in_1, msg_to_bit_it_13_vnu_83_in_2, msg_to_bit_it_13_vnu_84_in_0, msg_to_bit_it_13_vnu_84_in_1, msg_to_bit_it_13_vnu_84_in_2, msg_to_bit_it_13_vnu_85_in_0, msg_to_bit_it_13_vnu_85_in_1, msg_to_bit_it_13_vnu_85_in_2, msg_to_bit_it_13_vnu_86_in_0, msg_to_bit_it_13_vnu_86_in_1, msg_to_bit_it_13_vnu_86_in_2, msg_to_bit_it_13_vnu_87_in_0, msg_to_bit_it_13_vnu_87_in_1, msg_to_bit_it_13_vnu_87_in_2, msg_to_bit_it_13_vnu_88_in_0, msg_to_bit_it_13_vnu_88_in_1, msg_to_bit_it_13_vnu_88_in_2, msg_to_bit_it_13_vnu_89_in_0, msg_to_bit_it_13_vnu_89_in_1, msg_to_bit_it_13_vnu_89_in_2, msg_to_bit_it_13_vnu_90_in_0, msg_to_bit_it_13_vnu_90_in_1, msg_to_bit_it_13_vnu_90_in_2, msg_to_bit_it_13_vnu_91_in_0, msg_to_bit_it_13_vnu_91_in_1, msg_to_bit_it_13_vnu_91_in_2, msg_to_bit_it_13_vnu_92_in_0, msg_to_bit_it_13_vnu_92_in_1, msg_to_bit_it_13_vnu_92_in_2, msg_to_bit_it_13_vnu_93_in_0, msg_to_bit_it_13_vnu_93_in_1, msg_to_bit_it_13_vnu_93_in_2, msg_to_bit_it_13_vnu_94_in_0, msg_to_bit_it_13_vnu_94_in_1, msg_to_bit_it_13_vnu_94_in_2, msg_to_bit_it_13_vnu_95_in_0, msg_to_bit_it_13_vnu_95_in_1, msg_to_bit_it_13_vnu_95_in_2, msg_to_bit_it_13_vnu_96_in_0, msg_to_bit_it_13_vnu_96_in_1, msg_to_bit_it_13_vnu_96_in_2, msg_to_bit_it_13_vnu_97_in_0, msg_to_bit_it_13_vnu_97_in_1, msg_to_bit_it_13_vnu_97_in_2, msg_to_bit_it_13_vnu_98_in_0, msg_to_bit_it_13_vnu_98_in_1, msg_to_bit_it_13_vnu_98_in_2, msg_to_bit_it_13_vnu_99_in_0, msg_to_bit_it_13_vnu_99_in_1, msg_to_bit_it_13_vnu_99_in_2, msg_to_bit_it_13_vnu_100_in_0, msg_to_bit_it_13_vnu_100_in_1, msg_to_bit_it_13_vnu_100_in_2, msg_to_bit_it_13_vnu_101_in_0, msg_to_bit_it_13_vnu_101_in_1, msg_to_bit_it_13_vnu_101_in_2, msg_to_bit_it_13_vnu_102_in_0, msg_to_bit_it_13_vnu_102_in_1, msg_to_bit_it_13_vnu_102_in_2, msg_to_bit_it_13_vnu_103_in_0, msg_to_bit_it_13_vnu_103_in_1, msg_to_bit_it_13_vnu_103_in_2, msg_to_bit_it_13_vnu_104_in_0, msg_to_bit_it_13_vnu_104_in_1, msg_to_bit_it_13_vnu_104_in_2, msg_to_bit_it_13_vnu_105_in_0, msg_to_bit_it_13_vnu_105_in_1, msg_to_bit_it_13_vnu_105_in_2, msg_to_bit_it_13_vnu_106_in_0, msg_to_bit_it_13_vnu_106_in_1, msg_to_bit_it_13_vnu_106_in_2, msg_to_bit_it_13_vnu_107_in_0, msg_to_bit_it_13_vnu_107_in_1, msg_to_bit_it_13_vnu_107_in_2, msg_to_bit_it_13_vnu_108_in_0, msg_to_bit_it_13_vnu_108_in_1, msg_to_bit_it_13_vnu_108_in_2, msg_to_bit_it_13_vnu_109_in_0, msg_to_bit_it_13_vnu_109_in_1, msg_to_bit_it_13_vnu_109_in_2, msg_to_bit_it_13_vnu_110_in_0, msg_to_bit_it_13_vnu_110_in_1, msg_to_bit_it_13_vnu_110_in_2, msg_to_bit_it_13_vnu_111_in_0, msg_to_bit_it_13_vnu_111_in_1, msg_to_bit_it_13_vnu_111_in_2, msg_to_bit_it_13_vnu_112_in_0, msg_to_bit_it_13_vnu_112_in_1, msg_to_bit_it_13_vnu_112_in_2, msg_to_bit_it_13_vnu_113_in_0, msg_to_bit_it_13_vnu_113_in_1, msg_to_bit_it_13_vnu_113_in_2, msg_to_bit_it_13_vnu_114_in_0, msg_to_bit_it_13_vnu_114_in_1, msg_to_bit_it_13_vnu_114_in_2, msg_to_bit_it_13_vnu_115_in_0, msg_to_bit_it_13_vnu_115_in_1, msg_to_bit_it_13_vnu_115_in_2, msg_to_bit_it_13_vnu_116_in_0, msg_to_bit_it_13_vnu_116_in_1, msg_to_bit_it_13_vnu_116_in_2, msg_to_bit_it_13_vnu_117_in_0, msg_to_bit_it_13_vnu_117_in_1, msg_to_bit_it_13_vnu_117_in_2, msg_to_bit_it_13_vnu_118_in_0, msg_to_bit_it_13_vnu_118_in_1, msg_to_bit_it_13_vnu_118_in_2, msg_to_bit_it_13_vnu_119_in_0, msg_to_bit_it_13_vnu_119_in_1, msg_to_bit_it_13_vnu_119_in_2, msg_to_bit_it_13_vnu_120_in_0, msg_to_bit_it_13_vnu_120_in_1, msg_to_bit_it_13_vnu_120_in_2, msg_to_bit_it_13_vnu_121_in_0, msg_to_bit_it_13_vnu_121_in_1, msg_to_bit_it_13_vnu_121_in_2, msg_to_bit_it_13_vnu_122_in_0, msg_to_bit_it_13_vnu_122_in_1, msg_to_bit_it_13_vnu_122_in_2, msg_to_bit_it_13_vnu_123_in_0, msg_to_bit_it_13_vnu_123_in_1, msg_to_bit_it_13_vnu_123_in_2, msg_to_bit_it_13_vnu_124_in_0, msg_to_bit_it_13_vnu_124_in_1, msg_to_bit_it_13_vnu_124_in_2, msg_to_bit_it_13_vnu_125_in_0, msg_to_bit_it_13_vnu_125_in_1, msg_to_bit_it_13_vnu_125_in_2, msg_to_bit_it_13_vnu_126_in_0, msg_to_bit_it_13_vnu_126_in_1, msg_to_bit_it_13_vnu_126_in_2, msg_to_bit_it_13_vnu_127_in_0, msg_to_bit_it_13_vnu_127_in_1, msg_to_bit_it_13_vnu_127_in_2, msg_to_bit_it_13_vnu_128_in_0, msg_to_bit_it_13_vnu_128_in_1, msg_to_bit_it_13_vnu_128_in_2, msg_to_bit_it_13_vnu_129_in_0, msg_to_bit_it_13_vnu_129_in_1, msg_to_bit_it_13_vnu_129_in_2, msg_to_bit_it_13_vnu_130_in_0, msg_to_bit_it_13_vnu_130_in_1, msg_to_bit_it_13_vnu_130_in_2, msg_to_bit_it_13_vnu_131_in_0, msg_to_bit_it_13_vnu_131_in_1, msg_to_bit_it_13_vnu_131_in_2, msg_to_bit_it_13_vnu_132_in_0, msg_to_bit_it_13_vnu_132_in_1, msg_to_bit_it_13_vnu_132_in_2, msg_to_bit_it_13_vnu_133_in_0, msg_to_bit_it_13_vnu_133_in_1, msg_to_bit_it_13_vnu_133_in_2, msg_to_bit_it_13_vnu_134_in_0, msg_to_bit_it_13_vnu_134_in_1, msg_to_bit_it_13_vnu_134_in_2, msg_to_bit_it_13_vnu_135_in_0, msg_to_bit_it_13_vnu_135_in_1, msg_to_bit_it_13_vnu_135_in_2, msg_to_bit_it_13_vnu_136_in_0, msg_to_bit_it_13_vnu_136_in_1, msg_to_bit_it_13_vnu_136_in_2, msg_to_bit_it_13_vnu_137_in_0, msg_to_bit_it_13_vnu_137_in_1, msg_to_bit_it_13_vnu_137_in_2, msg_to_bit_it_13_vnu_138_in_0, msg_to_bit_it_13_vnu_138_in_1, msg_to_bit_it_13_vnu_138_in_2, msg_to_bit_it_13_vnu_139_in_0, msg_to_bit_it_13_vnu_139_in_1, msg_to_bit_it_13_vnu_139_in_2, msg_to_bit_it_13_vnu_140_in_0, msg_to_bit_it_13_vnu_140_in_1, msg_to_bit_it_13_vnu_140_in_2, msg_to_bit_it_13_vnu_141_in_0, msg_to_bit_it_13_vnu_141_in_1, msg_to_bit_it_13_vnu_141_in_2, msg_to_bit_it_13_vnu_142_in_0, msg_to_bit_it_13_vnu_142_in_1, msg_to_bit_it_13_vnu_142_in_2, msg_to_bit_it_13_vnu_143_in_0, msg_to_bit_it_13_vnu_143_in_1, msg_to_bit_it_13_vnu_143_in_2, msg_to_bit_it_13_vnu_144_in_0, msg_to_bit_it_13_vnu_144_in_1, msg_to_bit_it_13_vnu_144_in_2, msg_to_bit_it_13_vnu_145_in_0, msg_to_bit_it_13_vnu_145_in_1, msg_to_bit_it_13_vnu_145_in_2, msg_to_bit_it_13_vnu_146_in_0, msg_to_bit_it_13_vnu_146_in_1, msg_to_bit_it_13_vnu_146_in_2, msg_to_bit_it_13_vnu_147_in_0, msg_to_bit_it_13_vnu_147_in_1, msg_to_bit_it_13_vnu_147_in_2, msg_to_bit_it_13_vnu_148_in_0, msg_to_bit_it_13_vnu_148_in_1, msg_to_bit_it_13_vnu_148_in_2, msg_to_bit_it_13_vnu_149_in_0, msg_to_bit_it_13_vnu_149_in_1, msg_to_bit_it_13_vnu_149_in_2, msg_to_bit_it_13_vnu_150_in_0, msg_to_bit_it_13_vnu_150_in_1, msg_to_bit_it_13_vnu_150_in_2, msg_to_bit_it_13_vnu_151_in_0, msg_to_bit_it_13_vnu_151_in_1, msg_to_bit_it_13_vnu_151_in_2, msg_to_bit_it_13_vnu_152_in_0, msg_to_bit_it_13_vnu_152_in_1, msg_to_bit_it_13_vnu_152_in_2, msg_to_bit_it_13_vnu_153_in_0, msg_to_bit_it_13_vnu_153_in_1, msg_to_bit_it_13_vnu_153_in_2, msg_to_bit_it_13_vnu_154_in_0, msg_to_bit_it_13_vnu_154_in_1, msg_to_bit_it_13_vnu_154_in_2, msg_to_bit_it_13_vnu_155_in_0, msg_to_bit_it_13_vnu_155_in_1, msg_to_bit_it_13_vnu_155_in_2, msg_to_bit_it_13_vnu_156_in_0, msg_to_bit_it_13_vnu_156_in_1, msg_to_bit_it_13_vnu_156_in_2, msg_to_bit_it_13_vnu_157_in_0, msg_to_bit_it_13_vnu_157_in_1, msg_to_bit_it_13_vnu_157_in_2, msg_to_bit_it_13_vnu_158_in_0, msg_to_bit_it_13_vnu_158_in_1, msg_to_bit_it_13_vnu_158_in_2, msg_to_bit_it_13_vnu_159_in_0, msg_to_bit_it_13_vnu_159_in_1, msg_to_bit_it_13_vnu_159_in_2, msg_to_bit_it_13_vnu_160_in_0, msg_to_bit_it_13_vnu_160_in_1, msg_to_bit_it_13_vnu_160_in_2, msg_to_bit_it_13_vnu_161_in_0, msg_to_bit_it_13_vnu_161_in_1, msg_to_bit_it_13_vnu_161_in_2, msg_to_bit_it_13_vnu_162_in_0, msg_to_bit_it_13_vnu_162_in_1, msg_to_bit_it_13_vnu_162_in_2, msg_to_bit_it_13_vnu_163_in_0, msg_to_bit_it_13_vnu_163_in_1, msg_to_bit_it_13_vnu_163_in_2, msg_to_bit_it_13_vnu_164_in_0, msg_to_bit_it_13_vnu_164_in_1, msg_to_bit_it_13_vnu_164_in_2, msg_to_bit_it_13_vnu_165_in_0, msg_to_bit_it_13_vnu_165_in_1, msg_to_bit_it_13_vnu_165_in_2, msg_to_bit_it_13_vnu_166_in_0, msg_to_bit_it_13_vnu_166_in_1, msg_to_bit_it_13_vnu_166_in_2, msg_to_bit_it_13_vnu_167_in_0, msg_to_bit_it_13_vnu_167_in_1, msg_to_bit_it_13_vnu_167_in_2, msg_to_bit_it_13_vnu_168_in_0, msg_to_bit_it_13_vnu_168_in_1, msg_to_bit_it_13_vnu_168_in_2, msg_to_bit_it_13_vnu_169_in_0, msg_to_bit_it_13_vnu_169_in_1, msg_to_bit_it_13_vnu_169_in_2, msg_to_bit_it_13_vnu_170_in_0, msg_to_bit_it_13_vnu_170_in_1, msg_to_bit_it_13_vnu_170_in_2, msg_to_bit_it_13_vnu_171_in_0, msg_to_bit_it_13_vnu_171_in_1, msg_to_bit_it_13_vnu_171_in_2, msg_to_bit_it_13_vnu_172_in_0, msg_to_bit_it_13_vnu_172_in_1, msg_to_bit_it_13_vnu_172_in_2, msg_to_bit_it_13_vnu_173_in_0, msg_to_bit_it_13_vnu_173_in_1, msg_to_bit_it_13_vnu_173_in_2, msg_to_bit_it_13_vnu_174_in_0, msg_to_bit_it_13_vnu_174_in_1, msg_to_bit_it_13_vnu_174_in_2, msg_to_bit_it_13_vnu_175_in_0, msg_to_bit_it_13_vnu_175_in_1, msg_to_bit_it_13_vnu_175_in_2, msg_to_bit_it_13_vnu_176_in_0, msg_to_bit_it_13_vnu_176_in_1, msg_to_bit_it_13_vnu_176_in_2, msg_to_bit_it_13_vnu_177_in_0, msg_to_bit_it_13_vnu_177_in_1, msg_to_bit_it_13_vnu_177_in_2, msg_to_bit_it_13_vnu_178_in_0, msg_to_bit_it_13_vnu_178_in_1, msg_to_bit_it_13_vnu_178_in_2, msg_to_bit_it_13_vnu_179_in_0, msg_to_bit_it_13_vnu_179_in_1, msg_to_bit_it_13_vnu_179_in_2, msg_to_bit_it_13_vnu_180_in_0, msg_to_bit_it_13_vnu_180_in_1, msg_to_bit_it_13_vnu_180_in_2, msg_to_bit_it_13_vnu_181_in_0, msg_to_bit_it_13_vnu_181_in_1, msg_to_bit_it_13_vnu_181_in_2, msg_to_bit_it_13_vnu_182_in_0, msg_to_bit_it_13_vnu_182_in_1, msg_to_bit_it_13_vnu_182_in_2, msg_to_bit_it_13_vnu_183_in_0, msg_to_bit_it_13_vnu_183_in_1, msg_to_bit_it_13_vnu_183_in_2, msg_to_bit_it_13_vnu_184_in_0, msg_to_bit_it_13_vnu_184_in_1, msg_to_bit_it_13_vnu_184_in_2, msg_to_bit_it_13_vnu_185_in_0, msg_to_bit_it_13_vnu_185_in_1, msg_to_bit_it_13_vnu_185_in_2, msg_to_bit_it_13_vnu_186_in_0, msg_to_bit_it_13_vnu_186_in_1, msg_to_bit_it_13_vnu_186_in_2, msg_to_bit_it_13_vnu_187_in_0, msg_to_bit_it_13_vnu_187_in_1, msg_to_bit_it_13_vnu_187_in_2, msg_to_bit_it_13_vnu_188_in_0, msg_to_bit_it_13_vnu_188_in_1, msg_to_bit_it_13_vnu_188_in_2, msg_to_bit_it_13_vnu_189_in_0, msg_to_bit_it_13_vnu_189_in_1, msg_to_bit_it_13_vnu_189_in_2, msg_to_bit_it_13_vnu_190_in_0, msg_to_bit_it_13_vnu_190_in_1, msg_to_bit_it_13_vnu_190_in_2, msg_to_bit_it_13_vnu_191_in_0, msg_to_bit_it_13_vnu_191_in_1, msg_to_bit_it_13_vnu_191_in_2, msg_to_bit_it_13_vnu_192_in_0, msg_to_bit_it_13_vnu_192_in_1, msg_to_bit_it_13_vnu_192_in_2, msg_to_bit_it_13_vnu_193_in_0, msg_to_bit_it_13_vnu_193_in_1, msg_to_bit_it_13_vnu_193_in_2, msg_to_bit_it_13_vnu_194_in_0, msg_to_bit_it_13_vnu_194_in_1, msg_to_bit_it_13_vnu_194_in_2, msg_to_bit_it_13_vnu_195_in_0, msg_to_bit_it_13_vnu_195_in_1, msg_to_bit_it_13_vnu_195_in_2, msg_to_bit_it_13_vnu_196_in_0, msg_to_bit_it_13_vnu_196_in_1, msg_to_bit_it_13_vnu_196_in_2, msg_to_bit_it_13_vnu_197_in_0, msg_to_bit_it_13_vnu_197_in_1, msg_to_bit_it_13_vnu_197_in_2, msg_to_bit_it_14_vnu_0_in_0, msg_to_bit_it_14_vnu_0_in_1, msg_to_bit_it_14_vnu_0_in_2, msg_to_bit_it_14_vnu_1_in_0, msg_to_bit_it_14_vnu_1_in_1, msg_to_bit_it_14_vnu_1_in_2, msg_to_bit_it_14_vnu_2_in_0, msg_to_bit_it_14_vnu_2_in_1, msg_to_bit_it_14_vnu_2_in_2, msg_to_bit_it_14_vnu_3_in_0, msg_to_bit_it_14_vnu_3_in_1, msg_to_bit_it_14_vnu_3_in_2, msg_to_bit_it_14_vnu_4_in_0, msg_to_bit_it_14_vnu_4_in_1, msg_to_bit_it_14_vnu_4_in_2, msg_to_bit_it_14_vnu_5_in_0, msg_to_bit_it_14_vnu_5_in_1, msg_to_bit_it_14_vnu_5_in_2, msg_to_bit_it_14_vnu_6_in_0, msg_to_bit_it_14_vnu_6_in_1, msg_to_bit_it_14_vnu_6_in_2, msg_to_bit_it_14_vnu_7_in_0, msg_to_bit_it_14_vnu_7_in_1, msg_to_bit_it_14_vnu_7_in_2, msg_to_bit_it_14_vnu_8_in_0, msg_to_bit_it_14_vnu_8_in_1, msg_to_bit_it_14_vnu_8_in_2, msg_to_bit_it_14_vnu_9_in_0, msg_to_bit_it_14_vnu_9_in_1, msg_to_bit_it_14_vnu_9_in_2, msg_to_bit_it_14_vnu_10_in_0, msg_to_bit_it_14_vnu_10_in_1, msg_to_bit_it_14_vnu_10_in_2, msg_to_bit_it_14_vnu_11_in_0, msg_to_bit_it_14_vnu_11_in_1, msg_to_bit_it_14_vnu_11_in_2, msg_to_bit_it_14_vnu_12_in_0, msg_to_bit_it_14_vnu_12_in_1, msg_to_bit_it_14_vnu_12_in_2, msg_to_bit_it_14_vnu_13_in_0, msg_to_bit_it_14_vnu_13_in_1, msg_to_bit_it_14_vnu_13_in_2, msg_to_bit_it_14_vnu_14_in_0, msg_to_bit_it_14_vnu_14_in_1, msg_to_bit_it_14_vnu_14_in_2, msg_to_bit_it_14_vnu_15_in_0, msg_to_bit_it_14_vnu_15_in_1, msg_to_bit_it_14_vnu_15_in_2, msg_to_bit_it_14_vnu_16_in_0, msg_to_bit_it_14_vnu_16_in_1, msg_to_bit_it_14_vnu_16_in_2, msg_to_bit_it_14_vnu_17_in_0, msg_to_bit_it_14_vnu_17_in_1, msg_to_bit_it_14_vnu_17_in_2, msg_to_bit_it_14_vnu_18_in_0, msg_to_bit_it_14_vnu_18_in_1, msg_to_bit_it_14_vnu_18_in_2, msg_to_bit_it_14_vnu_19_in_0, msg_to_bit_it_14_vnu_19_in_1, msg_to_bit_it_14_vnu_19_in_2, msg_to_bit_it_14_vnu_20_in_0, msg_to_bit_it_14_vnu_20_in_1, msg_to_bit_it_14_vnu_20_in_2, msg_to_bit_it_14_vnu_21_in_0, msg_to_bit_it_14_vnu_21_in_1, msg_to_bit_it_14_vnu_21_in_2, msg_to_bit_it_14_vnu_22_in_0, msg_to_bit_it_14_vnu_22_in_1, msg_to_bit_it_14_vnu_22_in_2, msg_to_bit_it_14_vnu_23_in_0, msg_to_bit_it_14_vnu_23_in_1, msg_to_bit_it_14_vnu_23_in_2, msg_to_bit_it_14_vnu_24_in_0, msg_to_bit_it_14_vnu_24_in_1, msg_to_bit_it_14_vnu_24_in_2, msg_to_bit_it_14_vnu_25_in_0, msg_to_bit_it_14_vnu_25_in_1, msg_to_bit_it_14_vnu_25_in_2, msg_to_bit_it_14_vnu_26_in_0, msg_to_bit_it_14_vnu_26_in_1, msg_to_bit_it_14_vnu_26_in_2, msg_to_bit_it_14_vnu_27_in_0, msg_to_bit_it_14_vnu_27_in_1, msg_to_bit_it_14_vnu_27_in_2, msg_to_bit_it_14_vnu_28_in_0, msg_to_bit_it_14_vnu_28_in_1, msg_to_bit_it_14_vnu_28_in_2, msg_to_bit_it_14_vnu_29_in_0, msg_to_bit_it_14_vnu_29_in_1, msg_to_bit_it_14_vnu_29_in_2, msg_to_bit_it_14_vnu_30_in_0, msg_to_bit_it_14_vnu_30_in_1, msg_to_bit_it_14_vnu_30_in_2, msg_to_bit_it_14_vnu_31_in_0, msg_to_bit_it_14_vnu_31_in_1, msg_to_bit_it_14_vnu_31_in_2, msg_to_bit_it_14_vnu_32_in_0, msg_to_bit_it_14_vnu_32_in_1, msg_to_bit_it_14_vnu_32_in_2, msg_to_bit_it_14_vnu_33_in_0, msg_to_bit_it_14_vnu_33_in_1, msg_to_bit_it_14_vnu_33_in_2, msg_to_bit_it_14_vnu_34_in_0, msg_to_bit_it_14_vnu_34_in_1, msg_to_bit_it_14_vnu_34_in_2, msg_to_bit_it_14_vnu_35_in_0, msg_to_bit_it_14_vnu_35_in_1, msg_to_bit_it_14_vnu_35_in_2, msg_to_bit_it_14_vnu_36_in_0, msg_to_bit_it_14_vnu_36_in_1, msg_to_bit_it_14_vnu_36_in_2, msg_to_bit_it_14_vnu_37_in_0, msg_to_bit_it_14_vnu_37_in_1, msg_to_bit_it_14_vnu_37_in_2, msg_to_bit_it_14_vnu_38_in_0, msg_to_bit_it_14_vnu_38_in_1, msg_to_bit_it_14_vnu_38_in_2, msg_to_bit_it_14_vnu_39_in_0, msg_to_bit_it_14_vnu_39_in_1, msg_to_bit_it_14_vnu_39_in_2, msg_to_bit_it_14_vnu_40_in_0, msg_to_bit_it_14_vnu_40_in_1, msg_to_bit_it_14_vnu_40_in_2, msg_to_bit_it_14_vnu_41_in_0, msg_to_bit_it_14_vnu_41_in_1, msg_to_bit_it_14_vnu_41_in_2, msg_to_bit_it_14_vnu_42_in_0, msg_to_bit_it_14_vnu_42_in_1, msg_to_bit_it_14_vnu_42_in_2, msg_to_bit_it_14_vnu_43_in_0, msg_to_bit_it_14_vnu_43_in_1, msg_to_bit_it_14_vnu_43_in_2, msg_to_bit_it_14_vnu_44_in_0, msg_to_bit_it_14_vnu_44_in_1, msg_to_bit_it_14_vnu_44_in_2, msg_to_bit_it_14_vnu_45_in_0, msg_to_bit_it_14_vnu_45_in_1, msg_to_bit_it_14_vnu_45_in_2, msg_to_bit_it_14_vnu_46_in_0, msg_to_bit_it_14_vnu_46_in_1, msg_to_bit_it_14_vnu_46_in_2, msg_to_bit_it_14_vnu_47_in_0, msg_to_bit_it_14_vnu_47_in_1, msg_to_bit_it_14_vnu_47_in_2, msg_to_bit_it_14_vnu_48_in_0, msg_to_bit_it_14_vnu_48_in_1, msg_to_bit_it_14_vnu_48_in_2, msg_to_bit_it_14_vnu_49_in_0, msg_to_bit_it_14_vnu_49_in_1, msg_to_bit_it_14_vnu_49_in_2, msg_to_bit_it_14_vnu_50_in_0, msg_to_bit_it_14_vnu_50_in_1, msg_to_bit_it_14_vnu_50_in_2, msg_to_bit_it_14_vnu_51_in_0, msg_to_bit_it_14_vnu_51_in_1, msg_to_bit_it_14_vnu_51_in_2, msg_to_bit_it_14_vnu_52_in_0, msg_to_bit_it_14_vnu_52_in_1, msg_to_bit_it_14_vnu_52_in_2, msg_to_bit_it_14_vnu_53_in_0, msg_to_bit_it_14_vnu_53_in_1, msg_to_bit_it_14_vnu_53_in_2, msg_to_bit_it_14_vnu_54_in_0, msg_to_bit_it_14_vnu_54_in_1, msg_to_bit_it_14_vnu_54_in_2, msg_to_bit_it_14_vnu_55_in_0, msg_to_bit_it_14_vnu_55_in_1, msg_to_bit_it_14_vnu_55_in_2, msg_to_bit_it_14_vnu_56_in_0, msg_to_bit_it_14_vnu_56_in_1, msg_to_bit_it_14_vnu_56_in_2, msg_to_bit_it_14_vnu_57_in_0, msg_to_bit_it_14_vnu_57_in_1, msg_to_bit_it_14_vnu_57_in_2, msg_to_bit_it_14_vnu_58_in_0, msg_to_bit_it_14_vnu_58_in_1, msg_to_bit_it_14_vnu_58_in_2, msg_to_bit_it_14_vnu_59_in_0, msg_to_bit_it_14_vnu_59_in_1, msg_to_bit_it_14_vnu_59_in_2, msg_to_bit_it_14_vnu_60_in_0, msg_to_bit_it_14_vnu_60_in_1, msg_to_bit_it_14_vnu_60_in_2, msg_to_bit_it_14_vnu_61_in_0, msg_to_bit_it_14_vnu_61_in_1, msg_to_bit_it_14_vnu_61_in_2, msg_to_bit_it_14_vnu_62_in_0, msg_to_bit_it_14_vnu_62_in_1, msg_to_bit_it_14_vnu_62_in_2, msg_to_bit_it_14_vnu_63_in_0, msg_to_bit_it_14_vnu_63_in_1, msg_to_bit_it_14_vnu_63_in_2, msg_to_bit_it_14_vnu_64_in_0, msg_to_bit_it_14_vnu_64_in_1, msg_to_bit_it_14_vnu_64_in_2, msg_to_bit_it_14_vnu_65_in_0, msg_to_bit_it_14_vnu_65_in_1, msg_to_bit_it_14_vnu_65_in_2, msg_to_bit_it_14_vnu_66_in_0, msg_to_bit_it_14_vnu_66_in_1, msg_to_bit_it_14_vnu_66_in_2, msg_to_bit_it_14_vnu_67_in_0, msg_to_bit_it_14_vnu_67_in_1, msg_to_bit_it_14_vnu_67_in_2, msg_to_bit_it_14_vnu_68_in_0, msg_to_bit_it_14_vnu_68_in_1, msg_to_bit_it_14_vnu_68_in_2, msg_to_bit_it_14_vnu_69_in_0, msg_to_bit_it_14_vnu_69_in_1, msg_to_bit_it_14_vnu_69_in_2, msg_to_bit_it_14_vnu_70_in_0, msg_to_bit_it_14_vnu_70_in_1, msg_to_bit_it_14_vnu_70_in_2, msg_to_bit_it_14_vnu_71_in_0, msg_to_bit_it_14_vnu_71_in_1, msg_to_bit_it_14_vnu_71_in_2, msg_to_bit_it_14_vnu_72_in_0, msg_to_bit_it_14_vnu_72_in_1, msg_to_bit_it_14_vnu_72_in_2, msg_to_bit_it_14_vnu_73_in_0, msg_to_bit_it_14_vnu_73_in_1, msg_to_bit_it_14_vnu_73_in_2, msg_to_bit_it_14_vnu_74_in_0, msg_to_bit_it_14_vnu_74_in_1, msg_to_bit_it_14_vnu_74_in_2, msg_to_bit_it_14_vnu_75_in_0, msg_to_bit_it_14_vnu_75_in_1, msg_to_bit_it_14_vnu_75_in_2, msg_to_bit_it_14_vnu_76_in_0, msg_to_bit_it_14_vnu_76_in_1, msg_to_bit_it_14_vnu_76_in_2, msg_to_bit_it_14_vnu_77_in_0, msg_to_bit_it_14_vnu_77_in_1, msg_to_bit_it_14_vnu_77_in_2, msg_to_bit_it_14_vnu_78_in_0, msg_to_bit_it_14_vnu_78_in_1, msg_to_bit_it_14_vnu_78_in_2, msg_to_bit_it_14_vnu_79_in_0, msg_to_bit_it_14_vnu_79_in_1, msg_to_bit_it_14_vnu_79_in_2, msg_to_bit_it_14_vnu_80_in_0, msg_to_bit_it_14_vnu_80_in_1, msg_to_bit_it_14_vnu_80_in_2, msg_to_bit_it_14_vnu_81_in_0, msg_to_bit_it_14_vnu_81_in_1, msg_to_bit_it_14_vnu_81_in_2, msg_to_bit_it_14_vnu_82_in_0, msg_to_bit_it_14_vnu_82_in_1, msg_to_bit_it_14_vnu_82_in_2, msg_to_bit_it_14_vnu_83_in_0, msg_to_bit_it_14_vnu_83_in_1, msg_to_bit_it_14_vnu_83_in_2, msg_to_bit_it_14_vnu_84_in_0, msg_to_bit_it_14_vnu_84_in_1, msg_to_bit_it_14_vnu_84_in_2, msg_to_bit_it_14_vnu_85_in_0, msg_to_bit_it_14_vnu_85_in_1, msg_to_bit_it_14_vnu_85_in_2, msg_to_bit_it_14_vnu_86_in_0, msg_to_bit_it_14_vnu_86_in_1, msg_to_bit_it_14_vnu_86_in_2, msg_to_bit_it_14_vnu_87_in_0, msg_to_bit_it_14_vnu_87_in_1, msg_to_bit_it_14_vnu_87_in_2, msg_to_bit_it_14_vnu_88_in_0, msg_to_bit_it_14_vnu_88_in_1, msg_to_bit_it_14_vnu_88_in_2, msg_to_bit_it_14_vnu_89_in_0, msg_to_bit_it_14_vnu_89_in_1, msg_to_bit_it_14_vnu_89_in_2, msg_to_bit_it_14_vnu_90_in_0, msg_to_bit_it_14_vnu_90_in_1, msg_to_bit_it_14_vnu_90_in_2, msg_to_bit_it_14_vnu_91_in_0, msg_to_bit_it_14_vnu_91_in_1, msg_to_bit_it_14_vnu_91_in_2, msg_to_bit_it_14_vnu_92_in_0, msg_to_bit_it_14_vnu_92_in_1, msg_to_bit_it_14_vnu_92_in_2, msg_to_bit_it_14_vnu_93_in_0, msg_to_bit_it_14_vnu_93_in_1, msg_to_bit_it_14_vnu_93_in_2, msg_to_bit_it_14_vnu_94_in_0, msg_to_bit_it_14_vnu_94_in_1, msg_to_bit_it_14_vnu_94_in_2, msg_to_bit_it_14_vnu_95_in_0, msg_to_bit_it_14_vnu_95_in_1, msg_to_bit_it_14_vnu_95_in_2, msg_to_bit_it_14_vnu_96_in_0, msg_to_bit_it_14_vnu_96_in_1, msg_to_bit_it_14_vnu_96_in_2, msg_to_bit_it_14_vnu_97_in_0, msg_to_bit_it_14_vnu_97_in_1, msg_to_bit_it_14_vnu_97_in_2, msg_to_bit_it_14_vnu_98_in_0, msg_to_bit_it_14_vnu_98_in_1, msg_to_bit_it_14_vnu_98_in_2, msg_to_bit_it_14_vnu_99_in_0, msg_to_bit_it_14_vnu_99_in_1, msg_to_bit_it_14_vnu_99_in_2, msg_to_bit_it_14_vnu_100_in_0, msg_to_bit_it_14_vnu_100_in_1, msg_to_bit_it_14_vnu_100_in_2, msg_to_bit_it_14_vnu_101_in_0, msg_to_bit_it_14_vnu_101_in_1, msg_to_bit_it_14_vnu_101_in_2, msg_to_bit_it_14_vnu_102_in_0, msg_to_bit_it_14_vnu_102_in_1, msg_to_bit_it_14_vnu_102_in_2, msg_to_bit_it_14_vnu_103_in_0, msg_to_bit_it_14_vnu_103_in_1, msg_to_bit_it_14_vnu_103_in_2, msg_to_bit_it_14_vnu_104_in_0, msg_to_bit_it_14_vnu_104_in_1, msg_to_bit_it_14_vnu_104_in_2, msg_to_bit_it_14_vnu_105_in_0, msg_to_bit_it_14_vnu_105_in_1, msg_to_bit_it_14_vnu_105_in_2, msg_to_bit_it_14_vnu_106_in_0, msg_to_bit_it_14_vnu_106_in_1, msg_to_bit_it_14_vnu_106_in_2, msg_to_bit_it_14_vnu_107_in_0, msg_to_bit_it_14_vnu_107_in_1, msg_to_bit_it_14_vnu_107_in_2, msg_to_bit_it_14_vnu_108_in_0, msg_to_bit_it_14_vnu_108_in_1, msg_to_bit_it_14_vnu_108_in_2, msg_to_bit_it_14_vnu_109_in_0, msg_to_bit_it_14_vnu_109_in_1, msg_to_bit_it_14_vnu_109_in_2, msg_to_bit_it_14_vnu_110_in_0, msg_to_bit_it_14_vnu_110_in_1, msg_to_bit_it_14_vnu_110_in_2, msg_to_bit_it_14_vnu_111_in_0, msg_to_bit_it_14_vnu_111_in_1, msg_to_bit_it_14_vnu_111_in_2, msg_to_bit_it_14_vnu_112_in_0, msg_to_bit_it_14_vnu_112_in_1, msg_to_bit_it_14_vnu_112_in_2, msg_to_bit_it_14_vnu_113_in_0, msg_to_bit_it_14_vnu_113_in_1, msg_to_bit_it_14_vnu_113_in_2, msg_to_bit_it_14_vnu_114_in_0, msg_to_bit_it_14_vnu_114_in_1, msg_to_bit_it_14_vnu_114_in_2, msg_to_bit_it_14_vnu_115_in_0, msg_to_bit_it_14_vnu_115_in_1, msg_to_bit_it_14_vnu_115_in_2, msg_to_bit_it_14_vnu_116_in_0, msg_to_bit_it_14_vnu_116_in_1, msg_to_bit_it_14_vnu_116_in_2, msg_to_bit_it_14_vnu_117_in_0, msg_to_bit_it_14_vnu_117_in_1, msg_to_bit_it_14_vnu_117_in_2, msg_to_bit_it_14_vnu_118_in_0, msg_to_bit_it_14_vnu_118_in_1, msg_to_bit_it_14_vnu_118_in_2, msg_to_bit_it_14_vnu_119_in_0, msg_to_bit_it_14_vnu_119_in_1, msg_to_bit_it_14_vnu_119_in_2, msg_to_bit_it_14_vnu_120_in_0, msg_to_bit_it_14_vnu_120_in_1, msg_to_bit_it_14_vnu_120_in_2, msg_to_bit_it_14_vnu_121_in_0, msg_to_bit_it_14_vnu_121_in_1, msg_to_bit_it_14_vnu_121_in_2, msg_to_bit_it_14_vnu_122_in_0, msg_to_bit_it_14_vnu_122_in_1, msg_to_bit_it_14_vnu_122_in_2, msg_to_bit_it_14_vnu_123_in_0, msg_to_bit_it_14_vnu_123_in_1, msg_to_bit_it_14_vnu_123_in_2, msg_to_bit_it_14_vnu_124_in_0, msg_to_bit_it_14_vnu_124_in_1, msg_to_bit_it_14_vnu_124_in_2, msg_to_bit_it_14_vnu_125_in_0, msg_to_bit_it_14_vnu_125_in_1, msg_to_bit_it_14_vnu_125_in_2, msg_to_bit_it_14_vnu_126_in_0, msg_to_bit_it_14_vnu_126_in_1, msg_to_bit_it_14_vnu_126_in_2, msg_to_bit_it_14_vnu_127_in_0, msg_to_bit_it_14_vnu_127_in_1, msg_to_bit_it_14_vnu_127_in_2, msg_to_bit_it_14_vnu_128_in_0, msg_to_bit_it_14_vnu_128_in_1, msg_to_bit_it_14_vnu_128_in_2, msg_to_bit_it_14_vnu_129_in_0, msg_to_bit_it_14_vnu_129_in_1, msg_to_bit_it_14_vnu_129_in_2, msg_to_bit_it_14_vnu_130_in_0, msg_to_bit_it_14_vnu_130_in_1, msg_to_bit_it_14_vnu_130_in_2, msg_to_bit_it_14_vnu_131_in_0, msg_to_bit_it_14_vnu_131_in_1, msg_to_bit_it_14_vnu_131_in_2, msg_to_bit_it_14_vnu_132_in_0, msg_to_bit_it_14_vnu_132_in_1, msg_to_bit_it_14_vnu_132_in_2, msg_to_bit_it_14_vnu_133_in_0, msg_to_bit_it_14_vnu_133_in_1, msg_to_bit_it_14_vnu_133_in_2, msg_to_bit_it_14_vnu_134_in_0, msg_to_bit_it_14_vnu_134_in_1, msg_to_bit_it_14_vnu_134_in_2, msg_to_bit_it_14_vnu_135_in_0, msg_to_bit_it_14_vnu_135_in_1, msg_to_bit_it_14_vnu_135_in_2, msg_to_bit_it_14_vnu_136_in_0, msg_to_bit_it_14_vnu_136_in_1, msg_to_bit_it_14_vnu_136_in_2, msg_to_bit_it_14_vnu_137_in_0, msg_to_bit_it_14_vnu_137_in_1, msg_to_bit_it_14_vnu_137_in_2, msg_to_bit_it_14_vnu_138_in_0, msg_to_bit_it_14_vnu_138_in_1, msg_to_bit_it_14_vnu_138_in_2, msg_to_bit_it_14_vnu_139_in_0, msg_to_bit_it_14_vnu_139_in_1, msg_to_bit_it_14_vnu_139_in_2, msg_to_bit_it_14_vnu_140_in_0, msg_to_bit_it_14_vnu_140_in_1, msg_to_bit_it_14_vnu_140_in_2, msg_to_bit_it_14_vnu_141_in_0, msg_to_bit_it_14_vnu_141_in_1, msg_to_bit_it_14_vnu_141_in_2, msg_to_bit_it_14_vnu_142_in_0, msg_to_bit_it_14_vnu_142_in_1, msg_to_bit_it_14_vnu_142_in_2, msg_to_bit_it_14_vnu_143_in_0, msg_to_bit_it_14_vnu_143_in_1, msg_to_bit_it_14_vnu_143_in_2, msg_to_bit_it_14_vnu_144_in_0, msg_to_bit_it_14_vnu_144_in_1, msg_to_bit_it_14_vnu_144_in_2, msg_to_bit_it_14_vnu_145_in_0, msg_to_bit_it_14_vnu_145_in_1, msg_to_bit_it_14_vnu_145_in_2, msg_to_bit_it_14_vnu_146_in_0, msg_to_bit_it_14_vnu_146_in_1, msg_to_bit_it_14_vnu_146_in_2, msg_to_bit_it_14_vnu_147_in_0, msg_to_bit_it_14_vnu_147_in_1, msg_to_bit_it_14_vnu_147_in_2, msg_to_bit_it_14_vnu_148_in_0, msg_to_bit_it_14_vnu_148_in_1, msg_to_bit_it_14_vnu_148_in_2, msg_to_bit_it_14_vnu_149_in_0, msg_to_bit_it_14_vnu_149_in_1, msg_to_bit_it_14_vnu_149_in_2, msg_to_bit_it_14_vnu_150_in_0, msg_to_bit_it_14_vnu_150_in_1, msg_to_bit_it_14_vnu_150_in_2, msg_to_bit_it_14_vnu_151_in_0, msg_to_bit_it_14_vnu_151_in_1, msg_to_bit_it_14_vnu_151_in_2, msg_to_bit_it_14_vnu_152_in_0, msg_to_bit_it_14_vnu_152_in_1, msg_to_bit_it_14_vnu_152_in_2, msg_to_bit_it_14_vnu_153_in_0, msg_to_bit_it_14_vnu_153_in_1, msg_to_bit_it_14_vnu_153_in_2, msg_to_bit_it_14_vnu_154_in_0, msg_to_bit_it_14_vnu_154_in_1, msg_to_bit_it_14_vnu_154_in_2, msg_to_bit_it_14_vnu_155_in_0, msg_to_bit_it_14_vnu_155_in_1, msg_to_bit_it_14_vnu_155_in_2, msg_to_bit_it_14_vnu_156_in_0, msg_to_bit_it_14_vnu_156_in_1, msg_to_bit_it_14_vnu_156_in_2, msg_to_bit_it_14_vnu_157_in_0, msg_to_bit_it_14_vnu_157_in_1, msg_to_bit_it_14_vnu_157_in_2, msg_to_bit_it_14_vnu_158_in_0, msg_to_bit_it_14_vnu_158_in_1, msg_to_bit_it_14_vnu_158_in_2, msg_to_bit_it_14_vnu_159_in_0, msg_to_bit_it_14_vnu_159_in_1, msg_to_bit_it_14_vnu_159_in_2, msg_to_bit_it_14_vnu_160_in_0, msg_to_bit_it_14_vnu_160_in_1, msg_to_bit_it_14_vnu_160_in_2, msg_to_bit_it_14_vnu_161_in_0, msg_to_bit_it_14_vnu_161_in_1, msg_to_bit_it_14_vnu_161_in_2, msg_to_bit_it_14_vnu_162_in_0, msg_to_bit_it_14_vnu_162_in_1, msg_to_bit_it_14_vnu_162_in_2, msg_to_bit_it_14_vnu_163_in_0, msg_to_bit_it_14_vnu_163_in_1, msg_to_bit_it_14_vnu_163_in_2, msg_to_bit_it_14_vnu_164_in_0, msg_to_bit_it_14_vnu_164_in_1, msg_to_bit_it_14_vnu_164_in_2, msg_to_bit_it_14_vnu_165_in_0, msg_to_bit_it_14_vnu_165_in_1, msg_to_bit_it_14_vnu_165_in_2, msg_to_bit_it_14_vnu_166_in_0, msg_to_bit_it_14_vnu_166_in_1, msg_to_bit_it_14_vnu_166_in_2, msg_to_bit_it_14_vnu_167_in_0, msg_to_bit_it_14_vnu_167_in_1, msg_to_bit_it_14_vnu_167_in_2, msg_to_bit_it_14_vnu_168_in_0, msg_to_bit_it_14_vnu_168_in_1, msg_to_bit_it_14_vnu_168_in_2, msg_to_bit_it_14_vnu_169_in_0, msg_to_bit_it_14_vnu_169_in_1, msg_to_bit_it_14_vnu_169_in_2, msg_to_bit_it_14_vnu_170_in_0, msg_to_bit_it_14_vnu_170_in_1, msg_to_bit_it_14_vnu_170_in_2, msg_to_bit_it_14_vnu_171_in_0, msg_to_bit_it_14_vnu_171_in_1, msg_to_bit_it_14_vnu_171_in_2, msg_to_bit_it_14_vnu_172_in_0, msg_to_bit_it_14_vnu_172_in_1, msg_to_bit_it_14_vnu_172_in_2, msg_to_bit_it_14_vnu_173_in_0, msg_to_bit_it_14_vnu_173_in_1, msg_to_bit_it_14_vnu_173_in_2, msg_to_bit_it_14_vnu_174_in_0, msg_to_bit_it_14_vnu_174_in_1, msg_to_bit_it_14_vnu_174_in_2, msg_to_bit_it_14_vnu_175_in_0, msg_to_bit_it_14_vnu_175_in_1, msg_to_bit_it_14_vnu_175_in_2, msg_to_bit_it_14_vnu_176_in_0, msg_to_bit_it_14_vnu_176_in_1, msg_to_bit_it_14_vnu_176_in_2, msg_to_bit_it_14_vnu_177_in_0, msg_to_bit_it_14_vnu_177_in_1, msg_to_bit_it_14_vnu_177_in_2, msg_to_bit_it_14_vnu_178_in_0, msg_to_bit_it_14_vnu_178_in_1, msg_to_bit_it_14_vnu_178_in_2, msg_to_bit_it_14_vnu_179_in_0, msg_to_bit_it_14_vnu_179_in_1, msg_to_bit_it_14_vnu_179_in_2, msg_to_bit_it_14_vnu_180_in_0, msg_to_bit_it_14_vnu_180_in_1, msg_to_bit_it_14_vnu_180_in_2, msg_to_bit_it_14_vnu_181_in_0, msg_to_bit_it_14_vnu_181_in_1, msg_to_bit_it_14_vnu_181_in_2, msg_to_bit_it_14_vnu_182_in_0, msg_to_bit_it_14_vnu_182_in_1, msg_to_bit_it_14_vnu_182_in_2, msg_to_bit_it_14_vnu_183_in_0, msg_to_bit_it_14_vnu_183_in_1, msg_to_bit_it_14_vnu_183_in_2, msg_to_bit_it_14_vnu_184_in_0, msg_to_bit_it_14_vnu_184_in_1, msg_to_bit_it_14_vnu_184_in_2, msg_to_bit_it_14_vnu_185_in_0, msg_to_bit_it_14_vnu_185_in_1, msg_to_bit_it_14_vnu_185_in_2, msg_to_bit_it_14_vnu_186_in_0, msg_to_bit_it_14_vnu_186_in_1, msg_to_bit_it_14_vnu_186_in_2, msg_to_bit_it_14_vnu_187_in_0, msg_to_bit_it_14_vnu_187_in_1, msg_to_bit_it_14_vnu_187_in_2, msg_to_bit_it_14_vnu_188_in_0, msg_to_bit_it_14_vnu_188_in_1, msg_to_bit_it_14_vnu_188_in_2, msg_to_bit_it_14_vnu_189_in_0, msg_to_bit_it_14_vnu_189_in_1, msg_to_bit_it_14_vnu_189_in_2, msg_to_bit_it_14_vnu_190_in_0, msg_to_bit_it_14_vnu_190_in_1, msg_to_bit_it_14_vnu_190_in_2, msg_to_bit_it_14_vnu_191_in_0, msg_to_bit_it_14_vnu_191_in_1, msg_to_bit_it_14_vnu_191_in_2, msg_to_bit_it_14_vnu_192_in_0, msg_to_bit_it_14_vnu_192_in_1, msg_to_bit_it_14_vnu_192_in_2, msg_to_bit_it_14_vnu_193_in_0, msg_to_bit_it_14_vnu_193_in_1, msg_to_bit_it_14_vnu_193_in_2, msg_to_bit_it_14_vnu_194_in_0, msg_to_bit_it_14_vnu_194_in_1, msg_to_bit_it_14_vnu_194_in_2, msg_to_bit_it_14_vnu_195_in_0, msg_to_bit_it_14_vnu_195_in_1, msg_to_bit_it_14_vnu_195_in_2, msg_to_bit_it_14_vnu_196_in_0, msg_to_bit_it_14_vnu_196_in_1, msg_to_bit_it_14_vnu_196_in_2, msg_to_bit_it_14_vnu_197_in_0, msg_to_bit_it_14_vnu_197_in_1, msg_to_bit_it_14_vnu_197_in_2, msg_to_bit_it_15_vnu_0_in_0, msg_to_bit_it_15_vnu_0_in_1, msg_to_bit_it_15_vnu_0_in_2, msg_to_bit_it_15_vnu_1_in_0, msg_to_bit_it_15_vnu_1_in_1, msg_to_bit_it_15_vnu_1_in_2, msg_to_bit_it_15_vnu_2_in_0, msg_to_bit_it_15_vnu_2_in_1, msg_to_bit_it_15_vnu_2_in_2, msg_to_bit_it_15_vnu_3_in_0, msg_to_bit_it_15_vnu_3_in_1, msg_to_bit_it_15_vnu_3_in_2, msg_to_bit_it_15_vnu_4_in_0, msg_to_bit_it_15_vnu_4_in_1, msg_to_bit_it_15_vnu_4_in_2, msg_to_bit_it_15_vnu_5_in_0, msg_to_bit_it_15_vnu_5_in_1, msg_to_bit_it_15_vnu_5_in_2, msg_to_bit_it_15_vnu_6_in_0, msg_to_bit_it_15_vnu_6_in_1, msg_to_bit_it_15_vnu_6_in_2, msg_to_bit_it_15_vnu_7_in_0, msg_to_bit_it_15_vnu_7_in_1, msg_to_bit_it_15_vnu_7_in_2, msg_to_bit_it_15_vnu_8_in_0, msg_to_bit_it_15_vnu_8_in_1, msg_to_bit_it_15_vnu_8_in_2, msg_to_bit_it_15_vnu_9_in_0, msg_to_bit_it_15_vnu_9_in_1, msg_to_bit_it_15_vnu_9_in_2, msg_to_bit_it_15_vnu_10_in_0, msg_to_bit_it_15_vnu_10_in_1, msg_to_bit_it_15_vnu_10_in_2, msg_to_bit_it_15_vnu_11_in_0, msg_to_bit_it_15_vnu_11_in_1, msg_to_bit_it_15_vnu_11_in_2, msg_to_bit_it_15_vnu_12_in_0, msg_to_bit_it_15_vnu_12_in_1, msg_to_bit_it_15_vnu_12_in_2, msg_to_bit_it_15_vnu_13_in_0, msg_to_bit_it_15_vnu_13_in_1, msg_to_bit_it_15_vnu_13_in_2, msg_to_bit_it_15_vnu_14_in_0, msg_to_bit_it_15_vnu_14_in_1, msg_to_bit_it_15_vnu_14_in_2, msg_to_bit_it_15_vnu_15_in_0, msg_to_bit_it_15_vnu_15_in_1, msg_to_bit_it_15_vnu_15_in_2, msg_to_bit_it_15_vnu_16_in_0, msg_to_bit_it_15_vnu_16_in_1, msg_to_bit_it_15_vnu_16_in_2, msg_to_bit_it_15_vnu_17_in_0, msg_to_bit_it_15_vnu_17_in_1, msg_to_bit_it_15_vnu_17_in_2, msg_to_bit_it_15_vnu_18_in_0, msg_to_bit_it_15_vnu_18_in_1, msg_to_bit_it_15_vnu_18_in_2, msg_to_bit_it_15_vnu_19_in_0, msg_to_bit_it_15_vnu_19_in_1, msg_to_bit_it_15_vnu_19_in_2, msg_to_bit_it_15_vnu_20_in_0, msg_to_bit_it_15_vnu_20_in_1, msg_to_bit_it_15_vnu_20_in_2, msg_to_bit_it_15_vnu_21_in_0, msg_to_bit_it_15_vnu_21_in_1, msg_to_bit_it_15_vnu_21_in_2, msg_to_bit_it_15_vnu_22_in_0, msg_to_bit_it_15_vnu_22_in_1, msg_to_bit_it_15_vnu_22_in_2, msg_to_bit_it_15_vnu_23_in_0, msg_to_bit_it_15_vnu_23_in_1, msg_to_bit_it_15_vnu_23_in_2, msg_to_bit_it_15_vnu_24_in_0, msg_to_bit_it_15_vnu_24_in_1, msg_to_bit_it_15_vnu_24_in_2, msg_to_bit_it_15_vnu_25_in_0, msg_to_bit_it_15_vnu_25_in_1, msg_to_bit_it_15_vnu_25_in_2, msg_to_bit_it_15_vnu_26_in_0, msg_to_bit_it_15_vnu_26_in_1, msg_to_bit_it_15_vnu_26_in_2, msg_to_bit_it_15_vnu_27_in_0, msg_to_bit_it_15_vnu_27_in_1, msg_to_bit_it_15_vnu_27_in_2, msg_to_bit_it_15_vnu_28_in_0, msg_to_bit_it_15_vnu_28_in_1, msg_to_bit_it_15_vnu_28_in_2, msg_to_bit_it_15_vnu_29_in_0, msg_to_bit_it_15_vnu_29_in_1, msg_to_bit_it_15_vnu_29_in_2, msg_to_bit_it_15_vnu_30_in_0, msg_to_bit_it_15_vnu_30_in_1, msg_to_bit_it_15_vnu_30_in_2, msg_to_bit_it_15_vnu_31_in_0, msg_to_bit_it_15_vnu_31_in_1, msg_to_bit_it_15_vnu_31_in_2, msg_to_bit_it_15_vnu_32_in_0, msg_to_bit_it_15_vnu_32_in_1, msg_to_bit_it_15_vnu_32_in_2, msg_to_bit_it_15_vnu_33_in_0, msg_to_bit_it_15_vnu_33_in_1, msg_to_bit_it_15_vnu_33_in_2, msg_to_bit_it_15_vnu_34_in_0, msg_to_bit_it_15_vnu_34_in_1, msg_to_bit_it_15_vnu_34_in_2, msg_to_bit_it_15_vnu_35_in_0, msg_to_bit_it_15_vnu_35_in_1, msg_to_bit_it_15_vnu_35_in_2, msg_to_bit_it_15_vnu_36_in_0, msg_to_bit_it_15_vnu_36_in_1, msg_to_bit_it_15_vnu_36_in_2, msg_to_bit_it_15_vnu_37_in_0, msg_to_bit_it_15_vnu_37_in_1, msg_to_bit_it_15_vnu_37_in_2, msg_to_bit_it_15_vnu_38_in_0, msg_to_bit_it_15_vnu_38_in_1, msg_to_bit_it_15_vnu_38_in_2, msg_to_bit_it_15_vnu_39_in_0, msg_to_bit_it_15_vnu_39_in_1, msg_to_bit_it_15_vnu_39_in_2, msg_to_bit_it_15_vnu_40_in_0, msg_to_bit_it_15_vnu_40_in_1, msg_to_bit_it_15_vnu_40_in_2, msg_to_bit_it_15_vnu_41_in_0, msg_to_bit_it_15_vnu_41_in_1, msg_to_bit_it_15_vnu_41_in_2, msg_to_bit_it_15_vnu_42_in_0, msg_to_bit_it_15_vnu_42_in_1, msg_to_bit_it_15_vnu_42_in_2, msg_to_bit_it_15_vnu_43_in_0, msg_to_bit_it_15_vnu_43_in_1, msg_to_bit_it_15_vnu_43_in_2, msg_to_bit_it_15_vnu_44_in_0, msg_to_bit_it_15_vnu_44_in_1, msg_to_bit_it_15_vnu_44_in_2, msg_to_bit_it_15_vnu_45_in_0, msg_to_bit_it_15_vnu_45_in_1, msg_to_bit_it_15_vnu_45_in_2, msg_to_bit_it_15_vnu_46_in_0, msg_to_bit_it_15_vnu_46_in_1, msg_to_bit_it_15_vnu_46_in_2, msg_to_bit_it_15_vnu_47_in_0, msg_to_bit_it_15_vnu_47_in_1, msg_to_bit_it_15_vnu_47_in_2, msg_to_bit_it_15_vnu_48_in_0, msg_to_bit_it_15_vnu_48_in_1, msg_to_bit_it_15_vnu_48_in_2, msg_to_bit_it_15_vnu_49_in_0, msg_to_bit_it_15_vnu_49_in_1, msg_to_bit_it_15_vnu_49_in_2, msg_to_bit_it_15_vnu_50_in_0, msg_to_bit_it_15_vnu_50_in_1, msg_to_bit_it_15_vnu_50_in_2, msg_to_bit_it_15_vnu_51_in_0, msg_to_bit_it_15_vnu_51_in_1, msg_to_bit_it_15_vnu_51_in_2, msg_to_bit_it_15_vnu_52_in_0, msg_to_bit_it_15_vnu_52_in_1, msg_to_bit_it_15_vnu_52_in_2, msg_to_bit_it_15_vnu_53_in_0, msg_to_bit_it_15_vnu_53_in_1, msg_to_bit_it_15_vnu_53_in_2, msg_to_bit_it_15_vnu_54_in_0, msg_to_bit_it_15_vnu_54_in_1, msg_to_bit_it_15_vnu_54_in_2, msg_to_bit_it_15_vnu_55_in_0, msg_to_bit_it_15_vnu_55_in_1, msg_to_bit_it_15_vnu_55_in_2, msg_to_bit_it_15_vnu_56_in_0, msg_to_bit_it_15_vnu_56_in_1, msg_to_bit_it_15_vnu_56_in_2, msg_to_bit_it_15_vnu_57_in_0, msg_to_bit_it_15_vnu_57_in_1, msg_to_bit_it_15_vnu_57_in_2, msg_to_bit_it_15_vnu_58_in_0, msg_to_bit_it_15_vnu_58_in_1, msg_to_bit_it_15_vnu_58_in_2, msg_to_bit_it_15_vnu_59_in_0, msg_to_bit_it_15_vnu_59_in_1, msg_to_bit_it_15_vnu_59_in_2, msg_to_bit_it_15_vnu_60_in_0, msg_to_bit_it_15_vnu_60_in_1, msg_to_bit_it_15_vnu_60_in_2, msg_to_bit_it_15_vnu_61_in_0, msg_to_bit_it_15_vnu_61_in_1, msg_to_bit_it_15_vnu_61_in_2, msg_to_bit_it_15_vnu_62_in_0, msg_to_bit_it_15_vnu_62_in_1, msg_to_bit_it_15_vnu_62_in_2, msg_to_bit_it_15_vnu_63_in_0, msg_to_bit_it_15_vnu_63_in_1, msg_to_bit_it_15_vnu_63_in_2, msg_to_bit_it_15_vnu_64_in_0, msg_to_bit_it_15_vnu_64_in_1, msg_to_bit_it_15_vnu_64_in_2, msg_to_bit_it_15_vnu_65_in_0, msg_to_bit_it_15_vnu_65_in_1, msg_to_bit_it_15_vnu_65_in_2, msg_to_bit_it_15_vnu_66_in_0, msg_to_bit_it_15_vnu_66_in_1, msg_to_bit_it_15_vnu_66_in_2, msg_to_bit_it_15_vnu_67_in_0, msg_to_bit_it_15_vnu_67_in_1, msg_to_bit_it_15_vnu_67_in_2, msg_to_bit_it_15_vnu_68_in_0, msg_to_bit_it_15_vnu_68_in_1, msg_to_bit_it_15_vnu_68_in_2, msg_to_bit_it_15_vnu_69_in_0, msg_to_bit_it_15_vnu_69_in_1, msg_to_bit_it_15_vnu_69_in_2, msg_to_bit_it_15_vnu_70_in_0, msg_to_bit_it_15_vnu_70_in_1, msg_to_bit_it_15_vnu_70_in_2, msg_to_bit_it_15_vnu_71_in_0, msg_to_bit_it_15_vnu_71_in_1, msg_to_bit_it_15_vnu_71_in_2, msg_to_bit_it_15_vnu_72_in_0, msg_to_bit_it_15_vnu_72_in_1, msg_to_bit_it_15_vnu_72_in_2, msg_to_bit_it_15_vnu_73_in_0, msg_to_bit_it_15_vnu_73_in_1, msg_to_bit_it_15_vnu_73_in_2, msg_to_bit_it_15_vnu_74_in_0, msg_to_bit_it_15_vnu_74_in_1, msg_to_bit_it_15_vnu_74_in_2, msg_to_bit_it_15_vnu_75_in_0, msg_to_bit_it_15_vnu_75_in_1, msg_to_bit_it_15_vnu_75_in_2, msg_to_bit_it_15_vnu_76_in_0, msg_to_bit_it_15_vnu_76_in_1, msg_to_bit_it_15_vnu_76_in_2, msg_to_bit_it_15_vnu_77_in_0, msg_to_bit_it_15_vnu_77_in_1, msg_to_bit_it_15_vnu_77_in_2, msg_to_bit_it_15_vnu_78_in_0, msg_to_bit_it_15_vnu_78_in_1, msg_to_bit_it_15_vnu_78_in_2, msg_to_bit_it_15_vnu_79_in_0, msg_to_bit_it_15_vnu_79_in_1, msg_to_bit_it_15_vnu_79_in_2, msg_to_bit_it_15_vnu_80_in_0, msg_to_bit_it_15_vnu_80_in_1, msg_to_bit_it_15_vnu_80_in_2, msg_to_bit_it_15_vnu_81_in_0, msg_to_bit_it_15_vnu_81_in_1, msg_to_bit_it_15_vnu_81_in_2, msg_to_bit_it_15_vnu_82_in_0, msg_to_bit_it_15_vnu_82_in_1, msg_to_bit_it_15_vnu_82_in_2, msg_to_bit_it_15_vnu_83_in_0, msg_to_bit_it_15_vnu_83_in_1, msg_to_bit_it_15_vnu_83_in_2, msg_to_bit_it_15_vnu_84_in_0, msg_to_bit_it_15_vnu_84_in_1, msg_to_bit_it_15_vnu_84_in_2, msg_to_bit_it_15_vnu_85_in_0, msg_to_bit_it_15_vnu_85_in_1, msg_to_bit_it_15_vnu_85_in_2, msg_to_bit_it_15_vnu_86_in_0, msg_to_bit_it_15_vnu_86_in_1, msg_to_bit_it_15_vnu_86_in_2, msg_to_bit_it_15_vnu_87_in_0, msg_to_bit_it_15_vnu_87_in_1, msg_to_bit_it_15_vnu_87_in_2, msg_to_bit_it_15_vnu_88_in_0, msg_to_bit_it_15_vnu_88_in_1, msg_to_bit_it_15_vnu_88_in_2, msg_to_bit_it_15_vnu_89_in_0, msg_to_bit_it_15_vnu_89_in_1, msg_to_bit_it_15_vnu_89_in_2, msg_to_bit_it_15_vnu_90_in_0, msg_to_bit_it_15_vnu_90_in_1, msg_to_bit_it_15_vnu_90_in_2, msg_to_bit_it_15_vnu_91_in_0, msg_to_bit_it_15_vnu_91_in_1, msg_to_bit_it_15_vnu_91_in_2, msg_to_bit_it_15_vnu_92_in_0, msg_to_bit_it_15_vnu_92_in_1, msg_to_bit_it_15_vnu_92_in_2, msg_to_bit_it_15_vnu_93_in_0, msg_to_bit_it_15_vnu_93_in_1, msg_to_bit_it_15_vnu_93_in_2, msg_to_bit_it_15_vnu_94_in_0, msg_to_bit_it_15_vnu_94_in_1, msg_to_bit_it_15_vnu_94_in_2, msg_to_bit_it_15_vnu_95_in_0, msg_to_bit_it_15_vnu_95_in_1, msg_to_bit_it_15_vnu_95_in_2, msg_to_bit_it_15_vnu_96_in_0, msg_to_bit_it_15_vnu_96_in_1, msg_to_bit_it_15_vnu_96_in_2, msg_to_bit_it_15_vnu_97_in_0, msg_to_bit_it_15_vnu_97_in_1, msg_to_bit_it_15_vnu_97_in_2, msg_to_bit_it_15_vnu_98_in_0, msg_to_bit_it_15_vnu_98_in_1, msg_to_bit_it_15_vnu_98_in_2, msg_to_bit_it_15_vnu_99_in_0, msg_to_bit_it_15_vnu_99_in_1, msg_to_bit_it_15_vnu_99_in_2, msg_to_bit_it_15_vnu_100_in_0, msg_to_bit_it_15_vnu_100_in_1, msg_to_bit_it_15_vnu_100_in_2, msg_to_bit_it_15_vnu_101_in_0, msg_to_bit_it_15_vnu_101_in_1, msg_to_bit_it_15_vnu_101_in_2, msg_to_bit_it_15_vnu_102_in_0, msg_to_bit_it_15_vnu_102_in_1, msg_to_bit_it_15_vnu_102_in_2, msg_to_bit_it_15_vnu_103_in_0, msg_to_bit_it_15_vnu_103_in_1, msg_to_bit_it_15_vnu_103_in_2, msg_to_bit_it_15_vnu_104_in_0, msg_to_bit_it_15_vnu_104_in_1, msg_to_bit_it_15_vnu_104_in_2, msg_to_bit_it_15_vnu_105_in_0, msg_to_bit_it_15_vnu_105_in_1, msg_to_bit_it_15_vnu_105_in_2, msg_to_bit_it_15_vnu_106_in_0, msg_to_bit_it_15_vnu_106_in_1, msg_to_bit_it_15_vnu_106_in_2, msg_to_bit_it_15_vnu_107_in_0, msg_to_bit_it_15_vnu_107_in_1, msg_to_bit_it_15_vnu_107_in_2, msg_to_bit_it_15_vnu_108_in_0, msg_to_bit_it_15_vnu_108_in_1, msg_to_bit_it_15_vnu_108_in_2, msg_to_bit_it_15_vnu_109_in_0, msg_to_bit_it_15_vnu_109_in_1, msg_to_bit_it_15_vnu_109_in_2, msg_to_bit_it_15_vnu_110_in_0, msg_to_bit_it_15_vnu_110_in_1, msg_to_bit_it_15_vnu_110_in_2, msg_to_bit_it_15_vnu_111_in_0, msg_to_bit_it_15_vnu_111_in_1, msg_to_bit_it_15_vnu_111_in_2, msg_to_bit_it_15_vnu_112_in_0, msg_to_bit_it_15_vnu_112_in_1, msg_to_bit_it_15_vnu_112_in_2, msg_to_bit_it_15_vnu_113_in_0, msg_to_bit_it_15_vnu_113_in_1, msg_to_bit_it_15_vnu_113_in_2, msg_to_bit_it_15_vnu_114_in_0, msg_to_bit_it_15_vnu_114_in_1, msg_to_bit_it_15_vnu_114_in_2, msg_to_bit_it_15_vnu_115_in_0, msg_to_bit_it_15_vnu_115_in_1, msg_to_bit_it_15_vnu_115_in_2, msg_to_bit_it_15_vnu_116_in_0, msg_to_bit_it_15_vnu_116_in_1, msg_to_bit_it_15_vnu_116_in_2, msg_to_bit_it_15_vnu_117_in_0, msg_to_bit_it_15_vnu_117_in_1, msg_to_bit_it_15_vnu_117_in_2, msg_to_bit_it_15_vnu_118_in_0, msg_to_bit_it_15_vnu_118_in_1, msg_to_bit_it_15_vnu_118_in_2, msg_to_bit_it_15_vnu_119_in_0, msg_to_bit_it_15_vnu_119_in_1, msg_to_bit_it_15_vnu_119_in_2, msg_to_bit_it_15_vnu_120_in_0, msg_to_bit_it_15_vnu_120_in_1, msg_to_bit_it_15_vnu_120_in_2, msg_to_bit_it_15_vnu_121_in_0, msg_to_bit_it_15_vnu_121_in_1, msg_to_bit_it_15_vnu_121_in_2, msg_to_bit_it_15_vnu_122_in_0, msg_to_bit_it_15_vnu_122_in_1, msg_to_bit_it_15_vnu_122_in_2, msg_to_bit_it_15_vnu_123_in_0, msg_to_bit_it_15_vnu_123_in_1, msg_to_bit_it_15_vnu_123_in_2, msg_to_bit_it_15_vnu_124_in_0, msg_to_bit_it_15_vnu_124_in_1, msg_to_bit_it_15_vnu_124_in_2, msg_to_bit_it_15_vnu_125_in_0, msg_to_bit_it_15_vnu_125_in_1, msg_to_bit_it_15_vnu_125_in_2, msg_to_bit_it_15_vnu_126_in_0, msg_to_bit_it_15_vnu_126_in_1, msg_to_bit_it_15_vnu_126_in_2, msg_to_bit_it_15_vnu_127_in_0, msg_to_bit_it_15_vnu_127_in_1, msg_to_bit_it_15_vnu_127_in_2, msg_to_bit_it_15_vnu_128_in_0, msg_to_bit_it_15_vnu_128_in_1, msg_to_bit_it_15_vnu_128_in_2, msg_to_bit_it_15_vnu_129_in_0, msg_to_bit_it_15_vnu_129_in_1, msg_to_bit_it_15_vnu_129_in_2, msg_to_bit_it_15_vnu_130_in_0, msg_to_bit_it_15_vnu_130_in_1, msg_to_bit_it_15_vnu_130_in_2, msg_to_bit_it_15_vnu_131_in_0, msg_to_bit_it_15_vnu_131_in_1, msg_to_bit_it_15_vnu_131_in_2, msg_to_bit_it_15_vnu_132_in_0, msg_to_bit_it_15_vnu_132_in_1, msg_to_bit_it_15_vnu_132_in_2, msg_to_bit_it_15_vnu_133_in_0, msg_to_bit_it_15_vnu_133_in_1, msg_to_bit_it_15_vnu_133_in_2, msg_to_bit_it_15_vnu_134_in_0, msg_to_bit_it_15_vnu_134_in_1, msg_to_bit_it_15_vnu_134_in_2, msg_to_bit_it_15_vnu_135_in_0, msg_to_bit_it_15_vnu_135_in_1, msg_to_bit_it_15_vnu_135_in_2, msg_to_bit_it_15_vnu_136_in_0, msg_to_bit_it_15_vnu_136_in_1, msg_to_bit_it_15_vnu_136_in_2, msg_to_bit_it_15_vnu_137_in_0, msg_to_bit_it_15_vnu_137_in_1, msg_to_bit_it_15_vnu_137_in_2, msg_to_bit_it_15_vnu_138_in_0, msg_to_bit_it_15_vnu_138_in_1, msg_to_bit_it_15_vnu_138_in_2, msg_to_bit_it_15_vnu_139_in_0, msg_to_bit_it_15_vnu_139_in_1, msg_to_bit_it_15_vnu_139_in_2, msg_to_bit_it_15_vnu_140_in_0, msg_to_bit_it_15_vnu_140_in_1, msg_to_bit_it_15_vnu_140_in_2, msg_to_bit_it_15_vnu_141_in_0, msg_to_bit_it_15_vnu_141_in_1, msg_to_bit_it_15_vnu_141_in_2, msg_to_bit_it_15_vnu_142_in_0, msg_to_bit_it_15_vnu_142_in_1, msg_to_bit_it_15_vnu_142_in_2, msg_to_bit_it_15_vnu_143_in_0, msg_to_bit_it_15_vnu_143_in_1, msg_to_bit_it_15_vnu_143_in_2, msg_to_bit_it_15_vnu_144_in_0, msg_to_bit_it_15_vnu_144_in_1, msg_to_bit_it_15_vnu_144_in_2, msg_to_bit_it_15_vnu_145_in_0, msg_to_bit_it_15_vnu_145_in_1, msg_to_bit_it_15_vnu_145_in_2, msg_to_bit_it_15_vnu_146_in_0, msg_to_bit_it_15_vnu_146_in_1, msg_to_bit_it_15_vnu_146_in_2, msg_to_bit_it_15_vnu_147_in_0, msg_to_bit_it_15_vnu_147_in_1, msg_to_bit_it_15_vnu_147_in_2, msg_to_bit_it_15_vnu_148_in_0, msg_to_bit_it_15_vnu_148_in_1, msg_to_bit_it_15_vnu_148_in_2, msg_to_bit_it_15_vnu_149_in_0, msg_to_bit_it_15_vnu_149_in_1, msg_to_bit_it_15_vnu_149_in_2, msg_to_bit_it_15_vnu_150_in_0, msg_to_bit_it_15_vnu_150_in_1, msg_to_bit_it_15_vnu_150_in_2, msg_to_bit_it_15_vnu_151_in_0, msg_to_bit_it_15_vnu_151_in_1, msg_to_bit_it_15_vnu_151_in_2, msg_to_bit_it_15_vnu_152_in_0, msg_to_bit_it_15_vnu_152_in_1, msg_to_bit_it_15_vnu_152_in_2, msg_to_bit_it_15_vnu_153_in_0, msg_to_bit_it_15_vnu_153_in_1, msg_to_bit_it_15_vnu_153_in_2, msg_to_bit_it_15_vnu_154_in_0, msg_to_bit_it_15_vnu_154_in_1, msg_to_bit_it_15_vnu_154_in_2, msg_to_bit_it_15_vnu_155_in_0, msg_to_bit_it_15_vnu_155_in_1, msg_to_bit_it_15_vnu_155_in_2, msg_to_bit_it_15_vnu_156_in_0, msg_to_bit_it_15_vnu_156_in_1, msg_to_bit_it_15_vnu_156_in_2, msg_to_bit_it_15_vnu_157_in_0, msg_to_bit_it_15_vnu_157_in_1, msg_to_bit_it_15_vnu_157_in_2, msg_to_bit_it_15_vnu_158_in_0, msg_to_bit_it_15_vnu_158_in_1, msg_to_bit_it_15_vnu_158_in_2, msg_to_bit_it_15_vnu_159_in_0, msg_to_bit_it_15_vnu_159_in_1, msg_to_bit_it_15_vnu_159_in_2, msg_to_bit_it_15_vnu_160_in_0, msg_to_bit_it_15_vnu_160_in_1, msg_to_bit_it_15_vnu_160_in_2, msg_to_bit_it_15_vnu_161_in_0, msg_to_bit_it_15_vnu_161_in_1, msg_to_bit_it_15_vnu_161_in_2, msg_to_bit_it_15_vnu_162_in_0, msg_to_bit_it_15_vnu_162_in_1, msg_to_bit_it_15_vnu_162_in_2, msg_to_bit_it_15_vnu_163_in_0, msg_to_bit_it_15_vnu_163_in_1, msg_to_bit_it_15_vnu_163_in_2, msg_to_bit_it_15_vnu_164_in_0, msg_to_bit_it_15_vnu_164_in_1, msg_to_bit_it_15_vnu_164_in_2, msg_to_bit_it_15_vnu_165_in_0, msg_to_bit_it_15_vnu_165_in_1, msg_to_bit_it_15_vnu_165_in_2, msg_to_bit_it_15_vnu_166_in_0, msg_to_bit_it_15_vnu_166_in_1, msg_to_bit_it_15_vnu_166_in_2, msg_to_bit_it_15_vnu_167_in_0, msg_to_bit_it_15_vnu_167_in_1, msg_to_bit_it_15_vnu_167_in_2, msg_to_bit_it_15_vnu_168_in_0, msg_to_bit_it_15_vnu_168_in_1, msg_to_bit_it_15_vnu_168_in_2, msg_to_bit_it_15_vnu_169_in_0, msg_to_bit_it_15_vnu_169_in_1, msg_to_bit_it_15_vnu_169_in_2, msg_to_bit_it_15_vnu_170_in_0, msg_to_bit_it_15_vnu_170_in_1, msg_to_bit_it_15_vnu_170_in_2, msg_to_bit_it_15_vnu_171_in_0, msg_to_bit_it_15_vnu_171_in_1, msg_to_bit_it_15_vnu_171_in_2, msg_to_bit_it_15_vnu_172_in_0, msg_to_bit_it_15_vnu_172_in_1, msg_to_bit_it_15_vnu_172_in_2, msg_to_bit_it_15_vnu_173_in_0, msg_to_bit_it_15_vnu_173_in_1, msg_to_bit_it_15_vnu_173_in_2, msg_to_bit_it_15_vnu_174_in_0, msg_to_bit_it_15_vnu_174_in_1, msg_to_bit_it_15_vnu_174_in_2, msg_to_bit_it_15_vnu_175_in_0, msg_to_bit_it_15_vnu_175_in_1, msg_to_bit_it_15_vnu_175_in_2, msg_to_bit_it_15_vnu_176_in_0, msg_to_bit_it_15_vnu_176_in_1, msg_to_bit_it_15_vnu_176_in_2, msg_to_bit_it_15_vnu_177_in_0, msg_to_bit_it_15_vnu_177_in_1, msg_to_bit_it_15_vnu_177_in_2, msg_to_bit_it_15_vnu_178_in_0, msg_to_bit_it_15_vnu_178_in_1, msg_to_bit_it_15_vnu_178_in_2, msg_to_bit_it_15_vnu_179_in_0, msg_to_bit_it_15_vnu_179_in_1, msg_to_bit_it_15_vnu_179_in_2, msg_to_bit_it_15_vnu_180_in_0, msg_to_bit_it_15_vnu_180_in_1, msg_to_bit_it_15_vnu_180_in_2, msg_to_bit_it_15_vnu_181_in_0, msg_to_bit_it_15_vnu_181_in_1, msg_to_bit_it_15_vnu_181_in_2, msg_to_bit_it_15_vnu_182_in_0, msg_to_bit_it_15_vnu_182_in_1, msg_to_bit_it_15_vnu_182_in_2, msg_to_bit_it_15_vnu_183_in_0, msg_to_bit_it_15_vnu_183_in_1, msg_to_bit_it_15_vnu_183_in_2, msg_to_bit_it_15_vnu_184_in_0, msg_to_bit_it_15_vnu_184_in_1, msg_to_bit_it_15_vnu_184_in_2, msg_to_bit_it_15_vnu_185_in_0, msg_to_bit_it_15_vnu_185_in_1, msg_to_bit_it_15_vnu_185_in_2, msg_to_bit_it_15_vnu_186_in_0, msg_to_bit_it_15_vnu_186_in_1, msg_to_bit_it_15_vnu_186_in_2, msg_to_bit_it_15_vnu_187_in_0, msg_to_bit_it_15_vnu_187_in_1, msg_to_bit_it_15_vnu_187_in_2, msg_to_bit_it_15_vnu_188_in_0, msg_to_bit_it_15_vnu_188_in_1, msg_to_bit_it_15_vnu_188_in_2, msg_to_bit_it_15_vnu_189_in_0, msg_to_bit_it_15_vnu_189_in_1, msg_to_bit_it_15_vnu_189_in_2, msg_to_bit_it_15_vnu_190_in_0, msg_to_bit_it_15_vnu_190_in_1, msg_to_bit_it_15_vnu_190_in_2, msg_to_bit_it_15_vnu_191_in_0, msg_to_bit_it_15_vnu_191_in_1, msg_to_bit_it_15_vnu_191_in_2, msg_to_bit_it_15_vnu_192_in_0, msg_to_bit_it_15_vnu_192_in_1, msg_to_bit_it_15_vnu_192_in_2, msg_to_bit_it_15_vnu_193_in_0, msg_to_bit_it_15_vnu_193_in_1, msg_to_bit_it_15_vnu_193_in_2, msg_to_bit_it_15_vnu_194_in_0, msg_to_bit_it_15_vnu_194_in_1, msg_to_bit_it_15_vnu_194_in_2, msg_to_bit_it_15_vnu_195_in_0, msg_to_bit_it_15_vnu_195_in_1, msg_to_bit_it_15_vnu_195_in_2, msg_to_bit_it_15_vnu_196_in_0, msg_to_bit_it_15_vnu_196_in_1, msg_to_bit_it_15_vnu_196_in_2, msg_to_bit_it_15_vnu_197_in_0, msg_to_bit_it_15_vnu_197_in_1, msg_to_bit_it_15_vnu_197_in_2, msg_to_bit_it_16_vnu_0_in_0, msg_to_bit_it_16_vnu_0_in_1, msg_to_bit_it_16_vnu_0_in_2, msg_to_bit_it_16_vnu_1_in_0, msg_to_bit_it_16_vnu_1_in_1, msg_to_bit_it_16_vnu_1_in_2, msg_to_bit_it_16_vnu_2_in_0, msg_to_bit_it_16_vnu_2_in_1, msg_to_bit_it_16_vnu_2_in_2, msg_to_bit_it_16_vnu_3_in_0, msg_to_bit_it_16_vnu_3_in_1, msg_to_bit_it_16_vnu_3_in_2, msg_to_bit_it_16_vnu_4_in_0, msg_to_bit_it_16_vnu_4_in_1, msg_to_bit_it_16_vnu_4_in_2, msg_to_bit_it_16_vnu_5_in_0, msg_to_bit_it_16_vnu_5_in_1, msg_to_bit_it_16_vnu_5_in_2, msg_to_bit_it_16_vnu_6_in_0, msg_to_bit_it_16_vnu_6_in_1, msg_to_bit_it_16_vnu_6_in_2, msg_to_bit_it_16_vnu_7_in_0, msg_to_bit_it_16_vnu_7_in_1, msg_to_bit_it_16_vnu_7_in_2, msg_to_bit_it_16_vnu_8_in_0, msg_to_bit_it_16_vnu_8_in_1, msg_to_bit_it_16_vnu_8_in_2, msg_to_bit_it_16_vnu_9_in_0, msg_to_bit_it_16_vnu_9_in_1, msg_to_bit_it_16_vnu_9_in_2, msg_to_bit_it_16_vnu_10_in_0, msg_to_bit_it_16_vnu_10_in_1, msg_to_bit_it_16_vnu_10_in_2, msg_to_bit_it_16_vnu_11_in_0, msg_to_bit_it_16_vnu_11_in_1, msg_to_bit_it_16_vnu_11_in_2, msg_to_bit_it_16_vnu_12_in_0, msg_to_bit_it_16_vnu_12_in_1, msg_to_bit_it_16_vnu_12_in_2, msg_to_bit_it_16_vnu_13_in_0, msg_to_bit_it_16_vnu_13_in_1, msg_to_bit_it_16_vnu_13_in_2, msg_to_bit_it_16_vnu_14_in_0, msg_to_bit_it_16_vnu_14_in_1, msg_to_bit_it_16_vnu_14_in_2, msg_to_bit_it_16_vnu_15_in_0, msg_to_bit_it_16_vnu_15_in_1, msg_to_bit_it_16_vnu_15_in_2, msg_to_bit_it_16_vnu_16_in_0, msg_to_bit_it_16_vnu_16_in_1, msg_to_bit_it_16_vnu_16_in_2, msg_to_bit_it_16_vnu_17_in_0, msg_to_bit_it_16_vnu_17_in_1, msg_to_bit_it_16_vnu_17_in_2, msg_to_bit_it_16_vnu_18_in_0, msg_to_bit_it_16_vnu_18_in_1, msg_to_bit_it_16_vnu_18_in_2, msg_to_bit_it_16_vnu_19_in_0, msg_to_bit_it_16_vnu_19_in_1, msg_to_bit_it_16_vnu_19_in_2, msg_to_bit_it_16_vnu_20_in_0, msg_to_bit_it_16_vnu_20_in_1, msg_to_bit_it_16_vnu_20_in_2, msg_to_bit_it_16_vnu_21_in_0, msg_to_bit_it_16_vnu_21_in_1, msg_to_bit_it_16_vnu_21_in_2, msg_to_bit_it_16_vnu_22_in_0, msg_to_bit_it_16_vnu_22_in_1, msg_to_bit_it_16_vnu_22_in_2, msg_to_bit_it_16_vnu_23_in_0, msg_to_bit_it_16_vnu_23_in_1, msg_to_bit_it_16_vnu_23_in_2, msg_to_bit_it_16_vnu_24_in_0, msg_to_bit_it_16_vnu_24_in_1, msg_to_bit_it_16_vnu_24_in_2, msg_to_bit_it_16_vnu_25_in_0, msg_to_bit_it_16_vnu_25_in_1, msg_to_bit_it_16_vnu_25_in_2, msg_to_bit_it_16_vnu_26_in_0, msg_to_bit_it_16_vnu_26_in_1, msg_to_bit_it_16_vnu_26_in_2, msg_to_bit_it_16_vnu_27_in_0, msg_to_bit_it_16_vnu_27_in_1, msg_to_bit_it_16_vnu_27_in_2, msg_to_bit_it_16_vnu_28_in_0, msg_to_bit_it_16_vnu_28_in_1, msg_to_bit_it_16_vnu_28_in_2, msg_to_bit_it_16_vnu_29_in_0, msg_to_bit_it_16_vnu_29_in_1, msg_to_bit_it_16_vnu_29_in_2, msg_to_bit_it_16_vnu_30_in_0, msg_to_bit_it_16_vnu_30_in_1, msg_to_bit_it_16_vnu_30_in_2, msg_to_bit_it_16_vnu_31_in_0, msg_to_bit_it_16_vnu_31_in_1, msg_to_bit_it_16_vnu_31_in_2, msg_to_bit_it_16_vnu_32_in_0, msg_to_bit_it_16_vnu_32_in_1, msg_to_bit_it_16_vnu_32_in_2, msg_to_bit_it_16_vnu_33_in_0, msg_to_bit_it_16_vnu_33_in_1, msg_to_bit_it_16_vnu_33_in_2, msg_to_bit_it_16_vnu_34_in_0, msg_to_bit_it_16_vnu_34_in_1, msg_to_bit_it_16_vnu_34_in_2, msg_to_bit_it_16_vnu_35_in_0, msg_to_bit_it_16_vnu_35_in_1, msg_to_bit_it_16_vnu_35_in_2, msg_to_bit_it_16_vnu_36_in_0, msg_to_bit_it_16_vnu_36_in_1, msg_to_bit_it_16_vnu_36_in_2, msg_to_bit_it_16_vnu_37_in_0, msg_to_bit_it_16_vnu_37_in_1, msg_to_bit_it_16_vnu_37_in_2, msg_to_bit_it_16_vnu_38_in_0, msg_to_bit_it_16_vnu_38_in_1, msg_to_bit_it_16_vnu_38_in_2, msg_to_bit_it_16_vnu_39_in_0, msg_to_bit_it_16_vnu_39_in_1, msg_to_bit_it_16_vnu_39_in_2, msg_to_bit_it_16_vnu_40_in_0, msg_to_bit_it_16_vnu_40_in_1, msg_to_bit_it_16_vnu_40_in_2, msg_to_bit_it_16_vnu_41_in_0, msg_to_bit_it_16_vnu_41_in_1, msg_to_bit_it_16_vnu_41_in_2, msg_to_bit_it_16_vnu_42_in_0, msg_to_bit_it_16_vnu_42_in_1, msg_to_bit_it_16_vnu_42_in_2, msg_to_bit_it_16_vnu_43_in_0, msg_to_bit_it_16_vnu_43_in_1, msg_to_bit_it_16_vnu_43_in_2, msg_to_bit_it_16_vnu_44_in_0, msg_to_bit_it_16_vnu_44_in_1, msg_to_bit_it_16_vnu_44_in_2, msg_to_bit_it_16_vnu_45_in_0, msg_to_bit_it_16_vnu_45_in_1, msg_to_bit_it_16_vnu_45_in_2, msg_to_bit_it_16_vnu_46_in_0, msg_to_bit_it_16_vnu_46_in_1, msg_to_bit_it_16_vnu_46_in_2, msg_to_bit_it_16_vnu_47_in_0, msg_to_bit_it_16_vnu_47_in_1, msg_to_bit_it_16_vnu_47_in_2, msg_to_bit_it_16_vnu_48_in_0, msg_to_bit_it_16_vnu_48_in_1, msg_to_bit_it_16_vnu_48_in_2, msg_to_bit_it_16_vnu_49_in_0, msg_to_bit_it_16_vnu_49_in_1, msg_to_bit_it_16_vnu_49_in_2, msg_to_bit_it_16_vnu_50_in_0, msg_to_bit_it_16_vnu_50_in_1, msg_to_bit_it_16_vnu_50_in_2, msg_to_bit_it_16_vnu_51_in_0, msg_to_bit_it_16_vnu_51_in_1, msg_to_bit_it_16_vnu_51_in_2, msg_to_bit_it_16_vnu_52_in_0, msg_to_bit_it_16_vnu_52_in_1, msg_to_bit_it_16_vnu_52_in_2, msg_to_bit_it_16_vnu_53_in_0, msg_to_bit_it_16_vnu_53_in_1, msg_to_bit_it_16_vnu_53_in_2, msg_to_bit_it_16_vnu_54_in_0, msg_to_bit_it_16_vnu_54_in_1, msg_to_bit_it_16_vnu_54_in_2, msg_to_bit_it_16_vnu_55_in_0, msg_to_bit_it_16_vnu_55_in_1, msg_to_bit_it_16_vnu_55_in_2, msg_to_bit_it_16_vnu_56_in_0, msg_to_bit_it_16_vnu_56_in_1, msg_to_bit_it_16_vnu_56_in_2, msg_to_bit_it_16_vnu_57_in_0, msg_to_bit_it_16_vnu_57_in_1, msg_to_bit_it_16_vnu_57_in_2, msg_to_bit_it_16_vnu_58_in_0, msg_to_bit_it_16_vnu_58_in_1, msg_to_bit_it_16_vnu_58_in_2, msg_to_bit_it_16_vnu_59_in_0, msg_to_bit_it_16_vnu_59_in_1, msg_to_bit_it_16_vnu_59_in_2, msg_to_bit_it_16_vnu_60_in_0, msg_to_bit_it_16_vnu_60_in_1, msg_to_bit_it_16_vnu_60_in_2, msg_to_bit_it_16_vnu_61_in_0, msg_to_bit_it_16_vnu_61_in_1, msg_to_bit_it_16_vnu_61_in_2, msg_to_bit_it_16_vnu_62_in_0, msg_to_bit_it_16_vnu_62_in_1, msg_to_bit_it_16_vnu_62_in_2, msg_to_bit_it_16_vnu_63_in_0, msg_to_bit_it_16_vnu_63_in_1, msg_to_bit_it_16_vnu_63_in_2, msg_to_bit_it_16_vnu_64_in_0, msg_to_bit_it_16_vnu_64_in_1, msg_to_bit_it_16_vnu_64_in_2, msg_to_bit_it_16_vnu_65_in_0, msg_to_bit_it_16_vnu_65_in_1, msg_to_bit_it_16_vnu_65_in_2, msg_to_bit_it_16_vnu_66_in_0, msg_to_bit_it_16_vnu_66_in_1, msg_to_bit_it_16_vnu_66_in_2, msg_to_bit_it_16_vnu_67_in_0, msg_to_bit_it_16_vnu_67_in_1, msg_to_bit_it_16_vnu_67_in_2, msg_to_bit_it_16_vnu_68_in_0, msg_to_bit_it_16_vnu_68_in_1, msg_to_bit_it_16_vnu_68_in_2, msg_to_bit_it_16_vnu_69_in_0, msg_to_bit_it_16_vnu_69_in_1, msg_to_bit_it_16_vnu_69_in_2, msg_to_bit_it_16_vnu_70_in_0, msg_to_bit_it_16_vnu_70_in_1, msg_to_bit_it_16_vnu_70_in_2, msg_to_bit_it_16_vnu_71_in_0, msg_to_bit_it_16_vnu_71_in_1, msg_to_bit_it_16_vnu_71_in_2, msg_to_bit_it_16_vnu_72_in_0, msg_to_bit_it_16_vnu_72_in_1, msg_to_bit_it_16_vnu_72_in_2, msg_to_bit_it_16_vnu_73_in_0, msg_to_bit_it_16_vnu_73_in_1, msg_to_bit_it_16_vnu_73_in_2, msg_to_bit_it_16_vnu_74_in_0, msg_to_bit_it_16_vnu_74_in_1, msg_to_bit_it_16_vnu_74_in_2, msg_to_bit_it_16_vnu_75_in_0, msg_to_bit_it_16_vnu_75_in_1, msg_to_bit_it_16_vnu_75_in_2, msg_to_bit_it_16_vnu_76_in_0, msg_to_bit_it_16_vnu_76_in_1, msg_to_bit_it_16_vnu_76_in_2, msg_to_bit_it_16_vnu_77_in_0, msg_to_bit_it_16_vnu_77_in_1, msg_to_bit_it_16_vnu_77_in_2, msg_to_bit_it_16_vnu_78_in_0, msg_to_bit_it_16_vnu_78_in_1, msg_to_bit_it_16_vnu_78_in_2, msg_to_bit_it_16_vnu_79_in_0, msg_to_bit_it_16_vnu_79_in_1, msg_to_bit_it_16_vnu_79_in_2, msg_to_bit_it_16_vnu_80_in_0, msg_to_bit_it_16_vnu_80_in_1, msg_to_bit_it_16_vnu_80_in_2, msg_to_bit_it_16_vnu_81_in_0, msg_to_bit_it_16_vnu_81_in_1, msg_to_bit_it_16_vnu_81_in_2, msg_to_bit_it_16_vnu_82_in_0, msg_to_bit_it_16_vnu_82_in_1, msg_to_bit_it_16_vnu_82_in_2, msg_to_bit_it_16_vnu_83_in_0, msg_to_bit_it_16_vnu_83_in_1, msg_to_bit_it_16_vnu_83_in_2, msg_to_bit_it_16_vnu_84_in_0, msg_to_bit_it_16_vnu_84_in_1, msg_to_bit_it_16_vnu_84_in_2, msg_to_bit_it_16_vnu_85_in_0, msg_to_bit_it_16_vnu_85_in_1, msg_to_bit_it_16_vnu_85_in_2, msg_to_bit_it_16_vnu_86_in_0, msg_to_bit_it_16_vnu_86_in_1, msg_to_bit_it_16_vnu_86_in_2, msg_to_bit_it_16_vnu_87_in_0, msg_to_bit_it_16_vnu_87_in_1, msg_to_bit_it_16_vnu_87_in_2, msg_to_bit_it_16_vnu_88_in_0, msg_to_bit_it_16_vnu_88_in_1, msg_to_bit_it_16_vnu_88_in_2, msg_to_bit_it_16_vnu_89_in_0, msg_to_bit_it_16_vnu_89_in_1, msg_to_bit_it_16_vnu_89_in_2, msg_to_bit_it_16_vnu_90_in_0, msg_to_bit_it_16_vnu_90_in_1, msg_to_bit_it_16_vnu_90_in_2, msg_to_bit_it_16_vnu_91_in_0, msg_to_bit_it_16_vnu_91_in_1, msg_to_bit_it_16_vnu_91_in_2, msg_to_bit_it_16_vnu_92_in_0, msg_to_bit_it_16_vnu_92_in_1, msg_to_bit_it_16_vnu_92_in_2, msg_to_bit_it_16_vnu_93_in_0, msg_to_bit_it_16_vnu_93_in_1, msg_to_bit_it_16_vnu_93_in_2, msg_to_bit_it_16_vnu_94_in_0, msg_to_bit_it_16_vnu_94_in_1, msg_to_bit_it_16_vnu_94_in_2, msg_to_bit_it_16_vnu_95_in_0, msg_to_bit_it_16_vnu_95_in_1, msg_to_bit_it_16_vnu_95_in_2, msg_to_bit_it_16_vnu_96_in_0, msg_to_bit_it_16_vnu_96_in_1, msg_to_bit_it_16_vnu_96_in_2, msg_to_bit_it_16_vnu_97_in_0, msg_to_bit_it_16_vnu_97_in_1, msg_to_bit_it_16_vnu_97_in_2, msg_to_bit_it_16_vnu_98_in_0, msg_to_bit_it_16_vnu_98_in_1, msg_to_bit_it_16_vnu_98_in_2, msg_to_bit_it_16_vnu_99_in_0, msg_to_bit_it_16_vnu_99_in_1, msg_to_bit_it_16_vnu_99_in_2, msg_to_bit_it_16_vnu_100_in_0, msg_to_bit_it_16_vnu_100_in_1, msg_to_bit_it_16_vnu_100_in_2, msg_to_bit_it_16_vnu_101_in_0, msg_to_bit_it_16_vnu_101_in_1, msg_to_bit_it_16_vnu_101_in_2, msg_to_bit_it_16_vnu_102_in_0, msg_to_bit_it_16_vnu_102_in_1, msg_to_bit_it_16_vnu_102_in_2, msg_to_bit_it_16_vnu_103_in_0, msg_to_bit_it_16_vnu_103_in_1, msg_to_bit_it_16_vnu_103_in_2, msg_to_bit_it_16_vnu_104_in_0, msg_to_bit_it_16_vnu_104_in_1, msg_to_bit_it_16_vnu_104_in_2, msg_to_bit_it_16_vnu_105_in_0, msg_to_bit_it_16_vnu_105_in_1, msg_to_bit_it_16_vnu_105_in_2, msg_to_bit_it_16_vnu_106_in_0, msg_to_bit_it_16_vnu_106_in_1, msg_to_bit_it_16_vnu_106_in_2, msg_to_bit_it_16_vnu_107_in_0, msg_to_bit_it_16_vnu_107_in_1, msg_to_bit_it_16_vnu_107_in_2, msg_to_bit_it_16_vnu_108_in_0, msg_to_bit_it_16_vnu_108_in_1, msg_to_bit_it_16_vnu_108_in_2, msg_to_bit_it_16_vnu_109_in_0, msg_to_bit_it_16_vnu_109_in_1, msg_to_bit_it_16_vnu_109_in_2, msg_to_bit_it_16_vnu_110_in_0, msg_to_bit_it_16_vnu_110_in_1, msg_to_bit_it_16_vnu_110_in_2, msg_to_bit_it_16_vnu_111_in_0, msg_to_bit_it_16_vnu_111_in_1, msg_to_bit_it_16_vnu_111_in_2, msg_to_bit_it_16_vnu_112_in_0, msg_to_bit_it_16_vnu_112_in_1, msg_to_bit_it_16_vnu_112_in_2, msg_to_bit_it_16_vnu_113_in_0, msg_to_bit_it_16_vnu_113_in_1, msg_to_bit_it_16_vnu_113_in_2, msg_to_bit_it_16_vnu_114_in_0, msg_to_bit_it_16_vnu_114_in_1, msg_to_bit_it_16_vnu_114_in_2, msg_to_bit_it_16_vnu_115_in_0, msg_to_bit_it_16_vnu_115_in_1, msg_to_bit_it_16_vnu_115_in_2, msg_to_bit_it_16_vnu_116_in_0, msg_to_bit_it_16_vnu_116_in_1, msg_to_bit_it_16_vnu_116_in_2, msg_to_bit_it_16_vnu_117_in_0, msg_to_bit_it_16_vnu_117_in_1, msg_to_bit_it_16_vnu_117_in_2, msg_to_bit_it_16_vnu_118_in_0, msg_to_bit_it_16_vnu_118_in_1, msg_to_bit_it_16_vnu_118_in_2, msg_to_bit_it_16_vnu_119_in_0, msg_to_bit_it_16_vnu_119_in_1, msg_to_bit_it_16_vnu_119_in_2, msg_to_bit_it_16_vnu_120_in_0, msg_to_bit_it_16_vnu_120_in_1, msg_to_bit_it_16_vnu_120_in_2, msg_to_bit_it_16_vnu_121_in_0, msg_to_bit_it_16_vnu_121_in_1, msg_to_bit_it_16_vnu_121_in_2, msg_to_bit_it_16_vnu_122_in_0, msg_to_bit_it_16_vnu_122_in_1, msg_to_bit_it_16_vnu_122_in_2, msg_to_bit_it_16_vnu_123_in_0, msg_to_bit_it_16_vnu_123_in_1, msg_to_bit_it_16_vnu_123_in_2, msg_to_bit_it_16_vnu_124_in_0, msg_to_bit_it_16_vnu_124_in_1, msg_to_bit_it_16_vnu_124_in_2, msg_to_bit_it_16_vnu_125_in_0, msg_to_bit_it_16_vnu_125_in_1, msg_to_bit_it_16_vnu_125_in_2, msg_to_bit_it_16_vnu_126_in_0, msg_to_bit_it_16_vnu_126_in_1, msg_to_bit_it_16_vnu_126_in_2, msg_to_bit_it_16_vnu_127_in_0, msg_to_bit_it_16_vnu_127_in_1, msg_to_bit_it_16_vnu_127_in_2, msg_to_bit_it_16_vnu_128_in_0, msg_to_bit_it_16_vnu_128_in_1, msg_to_bit_it_16_vnu_128_in_2, msg_to_bit_it_16_vnu_129_in_0, msg_to_bit_it_16_vnu_129_in_1, msg_to_bit_it_16_vnu_129_in_2, msg_to_bit_it_16_vnu_130_in_0, msg_to_bit_it_16_vnu_130_in_1, msg_to_bit_it_16_vnu_130_in_2, msg_to_bit_it_16_vnu_131_in_0, msg_to_bit_it_16_vnu_131_in_1, msg_to_bit_it_16_vnu_131_in_2, msg_to_bit_it_16_vnu_132_in_0, msg_to_bit_it_16_vnu_132_in_1, msg_to_bit_it_16_vnu_132_in_2, msg_to_bit_it_16_vnu_133_in_0, msg_to_bit_it_16_vnu_133_in_1, msg_to_bit_it_16_vnu_133_in_2, msg_to_bit_it_16_vnu_134_in_0, msg_to_bit_it_16_vnu_134_in_1, msg_to_bit_it_16_vnu_134_in_2, msg_to_bit_it_16_vnu_135_in_0, msg_to_bit_it_16_vnu_135_in_1, msg_to_bit_it_16_vnu_135_in_2, msg_to_bit_it_16_vnu_136_in_0, msg_to_bit_it_16_vnu_136_in_1, msg_to_bit_it_16_vnu_136_in_2, msg_to_bit_it_16_vnu_137_in_0, msg_to_bit_it_16_vnu_137_in_1, msg_to_bit_it_16_vnu_137_in_2, msg_to_bit_it_16_vnu_138_in_0, msg_to_bit_it_16_vnu_138_in_1, msg_to_bit_it_16_vnu_138_in_2, msg_to_bit_it_16_vnu_139_in_0, msg_to_bit_it_16_vnu_139_in_1, msg_to_bit_it_16_vnu_139_in_2, msg_to_bit_it_16_vnu_140_in_0, msg_to_bit_it_16_vnu_140_in_1, msg_to_bit_it_16_vnu_140_in_2, msg_to_bit_it_16_vnu_141_in_0, msg_to_bit_it_16_vnu_141_in_1, msg_to_bit_it_16_vnu_141_in_2, msg_to_bit_it_16_vnu_142_in_0, msg_to_bit_it_16_vnu_142_in_1, msg_to_bit_it_16_vnu_142_in_2, msg_to_bit_it_16_vnu_143_in_0, msg_to_bit_it_16_vnu_143_in_1, msg_to_bit_it_16_vnu_143_in_2, msg_to_bit_it_16_vnu_144_in_0, msg_to_bit_it_16_vnu_144_in_1, msg_to_bit_it_16_vnu_144_in_2, msg_to_bit_it_16_vnu_145_in_0, msg_to_bit_it_16_vnu_145_in_1, msg_to_bit_it_16_vnu_145_in_2, msg_to_bit_it_16_vnu_146_in_0, msg_to_bit_it_16_vnu_146_in_1, msg_to_bit_it_16_vnu_146_in_2, msg_to_bit_it_16_vnu_147_in_0, msg_to_bit_it_16_vnu_147_in_1, msg_to_bit_it_16_vnu_147_in_2, msg_to_bit_it_16_vnu_148_in_0, msg_to_bit_it_16_vnu_148_in_1, msg_to_bit_it_16_vnu_148_in_2, msg_to_bit_it_16_vnu_149_in_0, msg_to_bit_it_16_vnu_149_in_1, msg_to_bit_it_16_vnu_149_in_2, msg_to_bit_it_16_vnu_150_in_0, msg_to_bit_it_16_vnu_150_in_1, msg_to_bit_it_16_vnu_150_in_2, msg_to_bit_it_16_vnu_151_in_0, msg_to_bit_it_16_vnu_151_in_1, msg_to_bit_it_16_vnu_151_in_2, msg_to_bit_it_16_vnu_152_in_0, msg_to_bit_it_16_vnu_152_in_1, msg_to_bit_it_16_vnu_152_in_2, msg_to_bit_it_16_vnu_153_in_0, msg_to_bit_it_16_vnu_153_in_1, msg_to_bit_it_16_vnu_153_in_2, msg_to_bit_it_16_vnu_154_in_0, msg_to_bit_it_16_vnu_154_in_1, msg_to_bit_it_16_vnu_154_in_2, msg_to_bit_it_16_vnu_155_in_0, msg_to_bit_it_16_vnu_155_in_1, msg_to_bit_it_16_vnu_155_in_2, msg_to_bit_it_16_vnu_156_in_0, msg_to_bit_it_16_vnu_156_in_1, msg_to_bit_it_16_vnu_156_in_2, msg_to_bit_it_16_vnu_157_in_0, msg_to_bit_it_16_vnu_157_in_1, msg_to_bit_it_16_vnu_157_in_2, msg_to_bit_it_16_vnu_158_in_0, msg_to_bit_it_16_vnu_158_in_1, msg_to_bit_it_16_vnu_158_in_2, msg_to_bit_it_16_vnu_159_in_0, msg_to_bit_it_16_vnu_159_in_1, msg_to_bit_it_16_vnu_159_in_2, msg_to_bit_it_16_vnu_160_in_0, msg_to_bit_it_16_vnu_160_in_1, msg_to_bit_it_16_vnu_160_in_2, msg_to_bit_it_16_vnu_161_in_0, msg_to_bit_it_16_vnu_161_in_1, msg_to_bit_it_16_vnu_161_in_2, msg_to_bit_it_16_vnu_162_in_0, msg_to_bit_it_16_vnu_162_in_1, msg_to_bit_it_16_vnu_162_in_2, msg_to_bit_it_16_vnu_163_in_0, msg_to_bit_it_16_vnu_163_in_1, msg_to_bit_it_16_vnu_163_in_2, msg_to_bit_it_16_vnu_164_in_0, msg_to_bit_it_16_vnu_164_in_1, msg_to_bit_it_16_vnu_164_in_2, msg_to_bit_it_16_vnu_165_in_0, msg_to_bit_it_16_vnu_165_in_1, msg_to_bit_it_16_vnu_165_in_2, msg_to_bit_it_16_vnu_166_in_0, msg_to_bit_it_16_vnu_166_in_1, msg_to_bit_it_16_vnu_166_in_2, msg_to_bit_it_16_vnu_167_in_0, msg_to_bit_it_16_vnu_167_in_1, msg_to_bit_it_16_vnu_167_in_2, msg_to_bit_it_16_vnu_168_in_0, msg_to_bit_it_16_vnu_168_in_1, msg_to_bit_it_16_vnu_168_in_2, msg_to_bit_it_16_vnu_169_in_0, msg_to_bit_it_16_vnu_169_in_1, msg_to_bit_it_16_vnu_169_in_2, msg_to_bit_it_16_vnu_170_in_0, msg_to_bit_it_16_vnu_170_in_1, msg_to_bit_it_16_vnu_170_in_2, msg_to_bit_it_16_vnu_171_in_0, msg_to_bit_it_16_vnu_171_in_1, msg_to_bit_it_16_vnu_171_in_2, msg_to_bit_it_16_vnu_172_in_0, msg_to_bit_it_16_vnu_172_in_1, msg_to_bit_it_16_vnu_172_in_2, msg_to_bit_it_16_vnu_173_in_0, msg_to_bit_it_16_vnu_173_in_1, msg_to_bit_it_16_vnu_173_in_2, msg_to_bit_it_16_vnu_174_in_0, msg_to_bit_it_16_vnu_174_in_1, msg_to_bit_it_16_vnu_174_in_2, msg_to_bit_it_16_vnu_175_in_0, msg_to_bit_it_16_vnu_175_in_1, msg_to_bit_it_16_vnu_175_in_2, msg_to_bit_it_16_vnu_176_in_0, msg_to_bit_it_16_vnu_176_in_1, msg_to_bit_it_16_vnu_176_in_2, msg_to_bit_it_16_vnu_177_in_0, msg_to_bit_it_16_vnu_177_in_1, msg_to_bit_it_16_vnu_177_in_2, msg_to_bit_it_16_vnu_178_in_0, msg_to_bit_it_16_vnu_178_in_1, msg_to_bit_it_16_vnu_178_in_2, msg_to_bit_it_16_vnu_179_in_0, msg_to_bit_it_16_vnu_179_in_1, msg_to_bit_it_16_vnu_179_in_2, msg_to_bit_it_16_vnu_180_in_0, msg_to_bit_it_16_vnu_180_in_1, msg_to_bit_it_16_vnu_180_in_2, msg_to_bit_it_16_vnu_181_in_0, msg_to_bit_it_16_vnu_181_in_1, msg_to_bit_it_16_vnu_181_in_2, msg_to_bit_it_16_vnu_182_in_0, msg_to_bit_it_16_vnu_182_in_1, msg_to_bit_it_16_vnu_182_in_2, msg_to_bit_it_16_vnu_183_in_0, msg_to_bit_it_16_vnu_183_in_1, msg_to_bit_it_16_vnu_183_in_2, msg_to_bit_it_16_vnu_184_in_0, msg_to_bit_it_16_vnu_184_in_1, msg_to_bit_it_16_vnu_184_in_2, msg_to_bit_it_16_vnu_185_in_0, msg_to_bit_it_16_vnu_185_in_1, msg_to_bit_it_16_vnu_185_in_2, msg_to_bit_it_16_vnu_186_in_0, msg_to_bit_it_16_vnu_186_in_1, msg_to_bit_it_16_vnu_186_in_2, msg_to_bit_it_16_vnu_187_in_0, msg_to_bit_it_16_vnu_187_in_1, msg_to_bit_it_16_vnu_187_in_2, msg_to_bit_it_16_vnu_188_in_0, msg_to_bit_it_16_vnu_188_in_1, msg_to_bit_it_16_vnu_188_in_2, msg_to_bit_it_16_vnu_189_in_0, msg_to_bit_it_16_vnu_189_in_1, msg_to_bit_it_16_vnu_189_in_2, msg_to_bit_it_16_vnu_190_in_0, msg_to_bit_it_16_vnu_190_in_1, msg_to_bit_it_16_vnu_190_in_2, msg_to_bit_it_16_vnu_191_in_0, msg_to_bit_it_16_vnu_191_in_1, msg_to_bit_it_16_vnu_191_in_2, msg_to_bit_it_16_vnu_192_in_0, msg_to_bit_it_16_vnu_192_in_1, msg_to_bit_it_16_vnu_192_in_2, msg_to_bit_it_16_vnu_193_in_0, msg_to_bit_it_16_vnu_193_in_1, msg_to_bit_it_16_vnu_193_in_2, msg_to_bit_it_16_vnu_194_in_0, msg_to_bit_it_16_vnu_194_in_1, msg_to_bit_it_16_vnu_194_in_2, msg_to_bit_it_16_vnu_195_in_0, msg_to_bit_it_16_vnu_195_in_1, msg_to_bit_it_16_vnu_195_in_2, msg_to_bit_it_16_vnu_196_in_0, msg_to_bit_it_16_vnu_196_in_1, msg_to_bit_it_16_vnu_196_in_2, msg_to_bit_it_16_vnu_197_in_0, msg_to_bit_it_16_vnu_197_in_1, msg_to_bit_it_16_vnu_197_in_2, msg_to_bit_it_17_vnu_0_in_0, msg_to_bit_it_17_vnu_0_in_1, msg_to_bit_it_17_vnu_0_in_2, msg_to_bit_it_17_vnu_1_in_0, msg_to_bit_it_17_vnu_1_in_1, msg_to_bit_it_17_vnu_1_in_2, msg_to_bit_it_17_vnu_2_in_0, msg_to_bit_it_17_vnu_2_in_1, msg_to_bit_it_17_vnu_2_in_2, msg_to_bit_it_17_vnu_3_in_0, msg_to_bit_it_17_vnu_3_in_1, msg_to_bit_it_17_vnu_3_in_2, msg_to_bit_it_17_vnu_4_in_0, msg_to_bit_it_17_vnu_4_in_1, msg_to_bit_it_17_vnu_4_in_2, msg_to_bit_it_17_vnu_5_in_0, msg_to_bit_it_17_vnu_5_in_1, msg_to_bit_it_17_vnu_5_in_2, msg_to_bit_it_17_vnu_6_in_0, msg_to_bit_it_17_vnu_6_in_1, msg_to_bit_it_17_vnu_6_in_2, msg_to_bit_it_17_vnu_7_in_0, msg_to_bit_it_17_vnu_7_in_1, msg_to_bit_it_17_vnu_7_in_2, msg_to_bit_it_17_vnu_8_in_0, msg_to_bit_it_17_vnu_8_in_1, msg_to_bit_it_17_vnu_8_in_2, msg_to_bit_it_17_vnu_9_in_0, msg_to_bit_it_17_vnu_9_in_1, msg_to_bit_it_17_vnu_9_in_2, msg_to_bit_it_17_vnu_10_in_0, msg_to_bit_it_17_vnu_10_in_1, msg_to_bit_it_17_vnu_10_in_2, msg_to_bit_it_17_vnu_11_in_0, msg_to_bit_it_17_vnu_11_in_1, msg_to_bit_it_17_vnu_11_in_2, msg_to_bit_it_17_vnu_12_in_0, msg_to_bit_it_17_vnu_12_in_1, msg_to_bit_it_17_vnu_12_in_2, msg_to_bit_it_17_vnu_13_in_0, msg_to_bit_it_17_vnu_13_in_1, msg_to_bit_it_17_vnu_13_in_2, msg_to_bit_it_17_vnu_14_in_0, msg_to_bit_it_17_vnu_14_in_1, msg_to_bit_it_17_vnu_14_in_2, msg_to_bit_it_17_vnu_15_in_0, msg_to_bit_it_17_vnu_15_in_1, msg_to_bit_it_17_vnu_15_in_2, msg_to_bit_it_17_vnu_16_in_0, msg_to_bit_it_17_vnu_16_in_1, msg_to_bit_it_17_vnu_16_in_2, msg_to_bit_it_17_vnu_17_in_0, msg_to_bit_it_17_vnu_17_in_1, msg_to_bit_it_17_vnu_17_in_2, msg_to_bit_it_17_vnu_18_in_0, msg_to_bit_it_17_vnu_18_in_1, msg_to_bit_it_17_vnu_18_in_2, msg_to_bit_it_17_vnu_19_in_0, msg_to_bit_it_17_vnu_19_in_1, msg_to_bit_it_17_vnu_19_in_2, msg_to_bit_it_17_vnu_20_in_0, msg_to_bit_it_17_vnu_20_in_1, msg_to_bit_it_17_vnu_20_in_2, msg_to_bit_it_17_vnu_21_in_0, msg_to_bit_it_17_vnu_21_in_1, msg_to_bit_it_17_vnu_21_in_2, msg_to_bit_it_17_vnu_22_in_0, msg_to_bit_it_17_vnu_22_in_1, msg_to_bit_it_17_vnu_22_in_2, msg_to_bit_it_17_vnu_23_in_0, msg_to_bit_it_17_vnu_23_in_1, msg_to_bit_it_17_vnu_23_in_2, msg_to_bit_it_17_vnu_24_in_0, msg_to_bit_it_17_vnu_24_in_1, msg_to_bit_it_17_vnu_24_in_2, msg_to_bit_it_17_vnu_25_in_0, msg_to_bit_it_17_vnu_25_in_1, msg_to_bit_it_17_vnu_25_in_2, msg_to_bit_it_17_vnu_26_in_0, msg_to_bit_it_17_vnu_26_in_1, msg_to_bit_it_17_vnu_26_in_2, msg_to_bit_it_17_vnu_27_in_0, msg_to_bit_it_17_vnu_27_in_1, msg_to_bit_it_17_vnu_27_in_2, msg_to_bit_it_17_vnu_28_in_0, msg_to_bit_it_17_vnu_28_in_1, msg_to_bit_it_17_vnu_28_in_2, msg_to_bit_it_17_vnu_29_in_0, msg_to_bit_it_17_vnu_29_in_1, msg_to_bit_it_17_vnu_29_in_2, msg_to_bit_it_17_vnu_30_in_0, msg_to_bit_it_17_vnu_30_in_1, msg_to_bit_it_17_vnu_30_in_2, msg_to_bit_it_17_vnu_31_in_0, msg_to_bit_it_17_vnu_31_in_1, msg_to_bit_it_17_vnu_31_in_2, msg_to_bit_it_17_vnu_32_in_0, msg_to_bit_it_17_vnu_32_in_1, msg_to_bit_it_17_vnu_32_in_2, msg_to_bit_it_17_vnu_33_in_0, msg_to_bit_it_17_vnu_33_in_1, msg_to_bit_it_17_vnu_33_in_2, msg_to_bit_it_17_vnu_34_in_0, msg_to_bit_it_17_vnu_34_in_1, msg_to_bit_it_17_vnu_34_in_2, msg_to_bit_it_17_vnu_35_in_0, msg_to_bit_it_17_vnu_35_in_1, msg_to_bit_it_17_vnu_35_in_2, msg_to_bit_it_17_vnu_36_in_0, msg_to_bit_it_17_vnu_36_in_1, msg_to_bit_it_17_vnu_36_in_2, msg_to_bit_it_17_vnu_37_in_0, msg_to_bit_it_17_vnu_37_in_1, msg_to_bit_it_17_vnu_37_in_2, msg_to_bit_it_17_vnu_38_in_0, msg_to_bit_it_17_vnu_38_in_1, msg_to_bit_it_17_vnu_38_in_2, msg_to_bit_it_17_vnu_39_in_0, msg_to_bit_it_17_vnu_39_in_1, msg_to_bit_it_17_vnu_39_in_2, msg_to_bit_it_17_vnu_40_in_0, msg_to_bit_it_17_vnu_40_in_1, msg_to_bit_it_17_vnu_40_in_2, msg_to_bit_it_17_vnu_41_in_0, msg_to_bit_it_17_vnu_41_in_1, msg_to_bit_it_17_vnu_41_in_2, msg_to_bit_it_17_vnu_42_in_0, msg_to_bit_it_17_vnu_42_in_1, msg_to_bit_it_17_vnu_42_in_2, msg_to_bit_it_17_vnu_43_in_0, msg_to_bit_it_17_vnu_43_in_1, msg_to_bit_it_17_vnu_43_in_2, msg_to_bit_it_17_vnu_44_in_0, msg_to_bit_it_17_vnu_44_in_1, msg_to_bit_it_17_vnu_44_in_2, msg_to_bit_it_17_vnu_45_in_0, msg_to_bit_it_17_vnu_45_in_1, msg_to_bit_it_17_vnu_45_in_2, msg_to_bit_it_17_vnu_46_in_0, msg_to_bit_it_17_vnu_46_in_1, msg_to_bit_it_17_vnu_46_in_2, msg_to_bit_it_17_vnu_47_in_0, msg_to_bit_it_17_vnu_47_in_1, msg_to_bit_it_17_vnu_47_in_2, msg_to_bit_it_17_vnu_48_in_0, msg_to_bit_it_17_vnu_48_in_1, msg_to_bit_it_17_vnu_48_in_2, msg_to_bit_it_17_vnu_49_in_0, msg_to_bit_it_17_vnu_49_in_1, msg_to_bit_it_17_vnu_49_in_2, msg_to_bit_it_17_vnu_50_in_0, msg_to_bit_it_17_vnu_50_in_1, msg_to_bit_it_17_vnu_50_in_2, msg_to_bit_it_17_vnu_51_in_0, msg_to_bit_it_17_vnu_51_in_1, msg_to_bit_it_17_vnu_51_in_2, msg_to_bit_it_17_vnu_52_in_0, msg_to_bit_it_17_vnu_52_in_1, msg_to_bit_it_17_vnu_52_in_2, msg_to_bit_it_17_vnu_53_in_0, msg_to_bit_it_17_vnu_53_in_1, msg_to_bit_it_17_vnu_53_in_2, msg_to_bit_it_17_vnu_54_in_0, msg_to_bit_it_17_vnu_54_in_1, msg_to_bit_it_17_vnu_54_in_2, msg_to_bit_it_17_vnu_55_in_0, msg_to_bit_it_17_vnu_55_in_1, msg_to_bit_it_17_vnu_55_in_2, msg_to_bit_it_17_vnu_56_in_0, msg_to_bit_it_17_vnu_56_in_1, msg_to_bit_it_17_vnu_56_in_2, msg_to_bit_it_17_vnu_57_in_0, msg_to_bit_it_17_vnu_57_in_1, msg_to_bit_it_17_vnu_57_in_2, msg_to_bit_it_17_vnu_58_in_0, msg_to_bit_it_17_vnu_58_in_1, msg_to_bit_it_17_vnu_58_in_2, msg_to_bit_it_17_vnu_59_in_0, msg_to_bit_it_17_vnu_59_in_1, msg_to_bit_it_17_vnu_59_in_2, msg_to_bit_it_17_vnu_60_in_0, msg_to_bit_it_17_vnu_60_in_1, msg_to_bit_it_17_vnu_60_in_2, msg_to_bit_it_17_vnu_61_in_0, msg_to_bit_it_17_vnu_61_in_1, msg_to_bit_it_17_vnu_61_in_2, msg_to_bit_it_17_vnu_62_in_0, msg_to_bit_it_17_vnu_62_in_1, msg_to_bit_it_17_vnu_62_in_2, msg_to_bit_it_17_vnu_63_in_0, msg_to_bit_it_17_vnu_63_in_1, msg_to_bit_it_17_vnu_63_in_2, msg_to_bit_it_17_vnu_64_in_0, msg_to_bit_it_17_vnu_64_in_1, msg_to_bit_it_17_vnu_64_in_2, msg_to_bit_it_17_vnu_65_in_0, msg_to_bit_it_17_vnu_65_in_1, msg_to_bit_it_17_vnu_65_in_2, msg_to_bit_it_17_vnu_66_in_0, msg_to_bit_it_17_vnu_66_in_1, msg_to_bit_it_17_vnu_66_in_2, msg_to_bit_it_17_vnu_67_in_0, msg_to_bit_it_17_vnu_67_in_1, msg_to_bit_it_17_vnu_67_in_2, msg_to_bit_it_17_vnu_68_in_0, msg_to_bit_it_17_vnu_68_in_1, msg_to_bit_it_17_vnu_68_in_2, msg_to_bit_it_17_vnu_69_in_0, msg_to_bit_it_17_vnu_69_in_1, msg_to_bit_it_17_vnu_69_in_2, msg_to_bit_it_17_vnu_70_in_0, msg_to_bit_it_17_vnu_70_in_1, msg_to_bit_it_17_vnu_70_in_2, msg_to_bit_it_17_vnu_71_in_0, msg_to_bit_it_17_vnu_71_in_1, msg_to_bit_it_17_vnu_71_in_2, msg_to_bit_it_17_vnu_72_in_0, msg_to_bit_it_17_vnu_72_in_1, msg_to_bit_it_17_vnu_72_in_2, msg_to_bit_it_17_vnu_73_in_0, msg_to_bit_it_17_vnu_73_in_1, msg_to_bit_it_17_vnu_73_in_2, msg_to_bit_it_17_vnu_74_in_0, msg_to_bit_it_17_vnu_74_in_1, msg_to_bit_it_17_vnu_74_in_2, msg_to_bit_it_17_vnu_75_in_0, msg_to_bit_it_17_vnu_75_in_1, msg_to_bit_it_17_vnu_75_in_2, msg_to_bit_it_17_vnu_76_in_0, msg_to_bit_it_17_vnu_76_in_1, msg_to_bit_it_17_vnu_76_in_2, msg_to_bit_it_17_vnu_77_in_0, msg_to_bit_it_17_vnu_77_in_1, msg_to_bit_it_17_vnu_77_in_2, msg_to_bit_it_17_vnu_78_in_0, msg_to_bit_it_17_vnu_78_in_1, msg_to_bit_it_17_vnu_78_in_2, msg_to_bit_it_17_vnu_79_in_0, msg_to_bit_it_17_vnu_79_in_1, msg_to_bit_it_17_vnu_79_in_2, msg_to_bit_it_17_vnu_80_in_0, msg_to_bit_it_17_vnu_80_in_1, msg_to_bit_it_17_vnu_80_in_2, msg_to_bit_it_17_vnu_81_in_0, msg_to_bit_it_17_vnu_81_in_1, msg_to_bit_it_17_vnu_81_in_2, msg_to_bit_it_17_vnu_82_in_0, msg_to_bit_it_17_vnu_82_in_1, msg_to_bit_it_17_vnu_82_in_2, msg_to_bit_it_17_vnu_83_in_0, msg_to_bit_it_17_vnu_83_in_1, msg_to_bit_it_17_vnu_83_in_2, msg_to_bit_it_17_vnu_84_in_0, msg_to_bit_it_17_vnu_84_in_1, msg_to_bit_it_17_vnu_84_in_2, msg_to_bit_it_17_vnu_85_in_0, msg_to_bit_it_17_vnu_85_in_1, msg_to_bit_it_17_vnu_85_in_2, msg_to_bit_it_17_vnu_86_in_0, msg_to_bit_it_17_vnu_86_in_1, msg_to_bit_it_17_vnu_86_in_2, msg_to_bit_it_17_vnu_87_in_0, msg_to_bit_it_17_vnu_87_in_1, msg_to_bit_it_17_vnu_87_in_2, msg_to_bit_it_17_vnu_88_in_0, msg_to_bit_it_17_vnu_88_in_1, msg_to_bit_it_17_vnu_88_in_2, msg_to_bit_it_17_vnu_89_in_0, msg_to_bit_it_17_vnu_89_in_1, msg_to_bit_it_17_vnu_89_in_2, msg_to_bit_it_17_vnu_90_in_0, msg_to_bit_it_17_vnu_90_in_1, msg_to_bit_it_17_vnu_90_in_2, msg_to_bit_it_17_vnu_91_in_0, msg_to_bit_it_17_vnu_91_in_1, msg_to_bit_it_17_vnu_91_in_2, msg_to_bit_it_17_vnu_92_in_0, msg_to_bit_it_17_vnu_92_in_1, msg_to_bit_it_17_vnu_92_in_2, msg_to_bit_it_17_vnu_93_in_0, msg_to_bit_it_17_vnu_93_in_1, msg_to_bit_it_17_vnu_93_in_2, msg_to_bit_it_17_vnu_94_in_0, msg_to_bit_it_17_vnu_94_in_1, msg_to_bit_it_17_vnu_94_in_2, msg_to_bit_it_17_vnu_95_in_0, msg_to_bit_it_17_vnu_95_in_1, msg_to_bit_it_17_vnu_95_in_2, msg_to_bit_it_17_vnu_96_in_0, msg_to_bit_it_17_vnu_96_in_1, msg_to_bit_it_17_vnu_96_in_2, msg_to_bit_it_17_vnu_97_in_0, msg_to_bit_it_17_vnu_97_in_1, msg_to_bit_it_17_vnu_97_in_2, msg_to_bit_it_17_vnu_98_in_0, msg_to_bit_it_17_vnu_98_in_1, msg_to_bit_it_17_vnu_98_in_2, msg_to_bit_it_17_vnu_99_in_0, msg_to_bit_it_17_vnu_99_in_1, msg_to_bit_it_17_vnu_99_in_2, msg_to_bit_it_17_vnu_100_in_0, msg_to_bit_it_17_vnu_100_in_1, msg_to_bit_it_17_vnu_100_in_2, msg_to_bit_it_17_vnu_101_in_0, msg_to_bit_it_17_vnu_101_in_1, msg_to_bit_it_17_vnu_101_in_2, msg_to_bit_it_17_vnu_102_in_0, msg_to_bit_it_17_vnu_102_in_1, msg_to_bit_it_17_vnu_102_in_2, msg_to_bit_it_17_vnu_103_in_0, msg_to_bit_it_17_vnu_103_in_1, msg_to_bit_it_17_vnu_103_in_2, msg_to_bit_it_17_vnu_104_in_0, msg_to_bit_it_17_vnu_104_in_1, msg_to_bit_it_17_vnu_104_in_2, msg_to_bit_it_17_vnu_105_in_0, msg_to_bit_it_17_vnu_105_in_1, msg_to_bit_it_17_vnu_105_in_2, msg_to_bit_it_17_vnu_106_in_0, msg_to_bit_it_17_vnu_106_in_1, msg_to_bit_it_17_vnu_106_in_2, msg_to_bit_it_17_vnu_107_in_0, msg_to_bit_it_17_vnu_107_in_1, msg_to_bit_it_17_vnu_107_in_2, msg_to_bit_it_17_vnu_108_in_0, msg_to_bit_it_17_vnu_108_in_1, msg_to_bit_it_17_vnu_108_in_2, msg_to_bit_it_17_vnu_109_in_0, msg_to_bit_it_17_vnu_109_in_1, msg_to_bit_it_17_vnu_109_in_2, msg_to_bit_it_17_vnu_110_in_0, msg_to_bit_it_17_vnu_110_in_1, msg_to_bit_it_17_vnu_110_in_2, msg_to_bit_it_17_vnu_111_in_0, msg_to_bit_it_17_vnu_111_in_1, msg_to_bit_it_17_vnu_111_in_2, msg_to_bit_it_17_vnu_112_in_0, msg_to_bit_it_17_vnu_112_in_1, msg_to_bit_it_17_vnu_112_in_2, msg_to_bit_it_17_vnu_113_in_0, msg_to_bit_it_17_vnu_113_in_1, msg_to_bit_it_17_vnu_113_in_2, msg_to_bit_it_17_vnu_114_in_0, msg_to_bit_it_17_vnu_114_in_1, msg_to_bit_it_17_vnu_114_in_2, msg_to_bit_it_17_vnu_115_in_0, msg_to_bit_it_17_vnu_115_in_1, msg_to_bit_it_17_vnu_115_in_2, msg_to_bit_it_17_vnu_116_in_0, msg_to_bit_it_17_vnu_116_in_1, msg_to_bit_it_17_vnu_116_in_2, msg_to_bit_it_17_vnu_117_in_0, msg_to_bit_it_17_vnu_117_in_1, msg_to_bit_it_17_vnu_117_in_2, msg_to_bit_it_17_vnu_118_in_0, msg_to_bit_it_17_vnu_118_in_1, msg_to_bit_it_17_vnu_118_in_2, msg_to_bit_it_17_vnu_119_in_0, msg_to_bit_it_17_vnu_119_in_1, msg_to_bit_it_17_vnu_119_in_2, msg_to_bit_it_17_vnu_120_in_0, msg_to_bit_it_17_vnu_120_in_1, msg_to_bit_it_17_vnu_120_in_2, msg_to_bit_it_17_vnu_121_in_0, msg_to_bit_it_17_vnu_121_in_1, msg_to_bit_it_17_vnu_121_in_2, msg_to_bit_it_17_vnu_122_in_0, msg_to_bit_it_17_vnu_122_in_1, msg_to_bit_it_17_vnu_122_in_2, msg_to_bit_it_17_vnu_123_in_0, msg_to_bit_it_17_vnu_123_in_1, msg_to_bit_it_17_vnu_123_in_2, msg_to_bit_it_17_vnu_124_in_0, msg_to_bit_it_17_vnu_124_in_1, msg_to_bit_it_17_vnu_124_in_2, msg_to_bit_it_17_vnu_125_in_0, msg_to_bit_it_17_vnu_125_in_1, msg_to_bit_it_17_vnu_125_in_2, msg_to_bit_it_17_vnu_126_in_0, msg_to_bit_it_17_vnu_126_in_1, msg_to_bit_it_17_vnu_126_in_2, msg_to_bit_it_17_vnu_127_in_0, msg_to_bit_it_17_vnu_127_in_1, msg_to_bit_it_17_vnu_127_in_2, msg_to_bit_it_17_vnu_128_in_0, msg_to_bit_it_17_vnu_128_in_1, msg_to_bit_it_17_vnu_128_in_2, msg_to_bit_it_17_vnu_129_in_0, msg_to_bit_it_17_vnu_129_in_1, msg_to_bit_it_17_vnu_129_in_2, msg_to_bit_it_17_vnu_130_in_0, msg_to_bit_it_17_vnu_130_in_1, msg_to_bit_it_17_vnu_130_in_2, msg_to_bit_it_17_vnu_131_in_0, msg_to_bit_it_17_vnu_131_in_1, msg_to_bit_it_17_vnu_131_in_2, msg_to_bit_it_17_vnu_132_in_0, msg_to_bit_it_17_vnu_132_in_1, msg_to_bit_it_17_vnu_132_in_2, msg_to_bit_it_17_vnu_133_in_0, msg_to_bit_it_17_vnu_133_in_1, msg_to_bit_it_17_vnu_133_in_2, msg_to_bit_it_17_vnu_134_in_0, msg_to_bit_it_17_vnu_134_in_1, msg_to_bit_it_17_vnu_134_in_2, msg_to_bit_it_17_vnu_135_in_0, msg_to_bit_it_17_vnu_135_in_1, msg_to_bit_it_17_vnu_135_in_2, msg_to_bit_it_17_vnu_136_in_0, msg_to_bit_it_17_vnu_136_in_1, msg_to_bit_it_17_vnu_136_in_2, msg_to_bit_it_17_vnu_137_in_0, msg_to_bit_it_17_vnu_137_in_1, msg_to_bit_it_17_vnu_137_in_2, msg_to_bit_it_17_vnu_138_in_0, msg_to_bit_it_17_vnu_138_in_1, msg_to_bit_it_17_vnu_138_in_2, msg_to_bit_it_17_vnu_139_in_0, msg_to_bit_it_17_vnu_139_in_1, msg_to_bit_it_17_vnu_139_in_2, msg_to_bit_it_17_vnu_140_in_0, msg_to_bit_it_17_vnu_140_in_1, msg_to_bit_it_17_vnu_140_in_2, msg_to_bit_it_17_vnu_141_in_0, msg_to_bit_it_17_vnu_141_in_1, msg_to_bit_it_17_vnu_141_in_2, msg_to_bit_it_17_vnu_142_in_0, msg_to_bit_it_17_vnu_142_in_1, msg_to_bit_it_17_vnu_142_in_2, msg_to_bit_it_17_vnu_143_in_0, msg_to_bit_it_17_vnu_143_in_1, msg_to_bit_it_17_vnu_143_in_2, msg_to_bit_it_17_vnu_144_in_0, msg_to_bit_it_17_vnu_144_in_1, msg_to_bit_it_17_vnu_144_in_2, msg_to_bit_it_17_vnu_145_in_0, msg_to_bit_it_17_vnu_145_in_1, msg_to_bit_it_17_vnu_145_in_2, msg_to_bit_it_17_vnu_146_in_0, msg_to_bit_it_17_vnu_146_in_1, msg_to_bit_it_17_vnu_146_in_2, msg_to_bit_it_17_vnu_147_in_0, msg_to_bit_it_17_vnu_147_in_1, msg_to_bit_it_17_vnu_147_in_2, msg_to_bit_it_17_vnu_148_in_0, msg_to_bit_it_17_vnu_148_in_1, msg_to_bit_it_17_vnu_148_in_2, msg_to_bit_it_17_vnu_149_in_0, msg_to_bit_it_17_vnu_149_in_1, msg_to_bit_it_17_vnu_149_in_2, msg_to_bit_it_17_vnu_150_in_0, msg_to_bit_it_17_vnu_150_in_1, msg_to_bit_it_17_vnu_150_in_2, msg_to_bit_it_17_vnu_151_in_0, msg_to_bit_it_17_vnu_151_in_1, msg_to_bit_it_17_vnu_151_in_2, msg_to_bit_it_17_vnu_152_in_0, msg_to_bit_it_17_vnu_152_in_1, msg_to_bit_it_17_vnu_152_in_2, msg_to_bit_it_17_vnu_153_in_0, msg_to_bit_it_17_vnu_153_in_1, msg_to_bit_it_17_vnu_153_in_2, msg_to_bit_it_17_vnu_154_in_0, msg_to_bit_it_17_vnu_154_in_1, msg_to_bit_it_17_vnu_154_in_2, msg_to_bit_it_17_vnu_155_in_0, msg_to_bit_it_17_vnu_155_in_1, msg_to_bit_it_17_vnu_155_in_2, msg_to_bit_it_17_vnu_156_in_0, msg_to_bit_it_17_vnu_156_in_1, msg_to_bit_it_17_vnu_156_in_2, msg_to_bit_it_17_vnu_157_in_0, msg_to_bit_it_17_vnu_157_in_1, msg_to_bit_it_17_vnu_157_in_2, msg_to_bit_it_17_vnu_158_in_0, msg_to_bit_it_17_vnu_158_in_1, msg_to_bit_it_17_vnu_158_in_2, msg_to_bit_it_17_vnu_159_in_0, msg_to_bit_it_17_vnu_159_in_1, msg_to_bit_it_17_vnu_159_in_2, msg_to_bit_it_17_vnu_160_in_0, msg_to_bit_it_17_vnu_160_in_1, msg_to_bit_it_17_vnu_160_in_2, msg_to_bit_it_17_vnu_161_in_0, msg_to_bit_it_17_vnu_161_in_1, msg_to_bit_it_17_vnu_161_in_2, msg_to_bit_it_17_vnu_162_in_0, msg_to_bit_it_17_vnu_162_in_1, msg_to_bit_it_17_vnu_162_in_2, msg_to_bit_it_17_vnu_163_in_0, msg_to_bit_it_17_vnu_163_in_1, msg_to_bit_it_17_vnu_163_in_2, msg_to_bit_it_17_vnu_164_in_0, msg_to_bit_it_17_vnu_164_in_1, msg_to_bit_it_17_vnu_164_in_2, msg_to_bit_it_17_vnu_165_in_0, msg_to_bit_it_17_vnu_165_in_1, msg_to_bit_it_17_vnu_165_in_2, msg_to_bit_it_17_vnu_166_in_0, msg_to_bit_it_17_vnu_166_in_1, msg_to_bit_it_17_vnu_166_in_2, msg_to_bit_it_17_vnu_167_in_0, msg_to_bit_it_17_vnu_167_in_1, msg_to_bit_it_17_vnu_167_in_2, msg_to_bit_it_17_vnu_168_in_0, msg_to_bit_it_17_vnu_168_in_1, msg_to_bit_it_17_vnu_168_in_2, msg_to_bit_it_17_vnu_169_in_0, msg_to_bit_it_17_vnu_169_in_1, msg_to_bit_it_17_vnu_169_in_2, msg_to_bit_it_17_vnu_170_in_0, msg_to_bit_it_17_vnu_170_in_1, msg_to_bit_it_17_vnu_170_in_2, msg_to_bit_it_17_vnu_171_in_0, msg_to_bit_it_17_vnu_171_in_1, msg_to_bit_it_17_vnu_171_in_2, msg_to_bit_it_17_vnu_172_in_0, msg_to_bit_it_17_vnu_172_in_1, msg_to_bit_it_17_vnu_172_in_2, msg_to_bit_it_17_vnu_173_in_0, msg_to_bit_it_17_vnu_173_in_1, msg_to_bit_it_17_vnu_173_in_2, msg_to_bit_it_17_vnu_174_in_0, msg_to_bit_it_17_vnu_174_in_1, msg_to_bit_it_17_vnu_174_in_2, msg_to_bit_it_17_vnu_175_in_0, msg_to_bit_it_17_vnu_175_in_1, msg_to_bit_it_17_vnu_175_in_2, msg_to_bit_it_17_vnu_176_in_0, msg_to_bit_it_17_vnu_176_in_1, msg_to_bit_it_17_vnu_176_in_2, msg_to_bit_it_17_vnu_177_in_0, msg_to_bit_it_17_vnu_177_in_1, msg_to_bit_it_17_vnu_177_in_2, msg_to_bit_it_17_vnu_178_in_0, msg_to_bit_it_17_vnu_178_in_1, msg_to_bit_it_17_vnu_178_in_2, msg_to_bit_it_17_vnu_179_in_0, msg_to_bit_it_17_vnu_179_in_1, msg_to_bit_it_17_vnu_179_in_2, msg_to_bit_it_17_vnu_180_in_0, msg_to_bit_it_17_vnu_180_in_1, msg_to_bit_it_17_vnu_180_in_2, msg_to_bit_it_17_vnu_181_in_0, msg_to_bit_it_17_vnu_181_in_1, msg_to_bit_it_17_vnu_181_in_2, msg_to_bit_it_17_vnu_182_in_0, msg_to_bit_it_17_vnu_182_in_1, msg_to_bit_it_17_vnu_182_in_2, msg_to_bit_it_17_vnu_183_in_0, msg_to_bit_it_17_vnu_183_in_1, msg_to_bit_it_17_vnu_183_in_2, msg_to_bit_it_17_vnu_184_in_0, msg_to_bit_it_17_vnu_184_in_1, msg_to_bit_it_17_vnu_184_in_2, msg_to_bit_it_17_vnu_185_in_0, msg_to_bit_it_17_vnu_185_in_1, msg_to_bit_it_17_vnu_185_in_2, msg_to_bit_it_17_vnu_186_in_0, msg_to_bit_it_17_vnu_186_in_1, msg_to_bit_it_17_vnu_186_in_2, msg_to_bit_it_17_vnu_187_in_0, msg_to_bit_it_17_vnu_187_in_1, msg_to_bit_it_17_vnu_187_in_2, msg_to_bit_it_17_vnu_188_in_0, msg_to_bit_it_17_vnu_188_in_1, msg_to_bit_it_17_vnu_188_in_2, msg_to_bit_it_17_vnu_189_in_0, msg_to_bit_it_17_vnu_189_in_1, msg_to_bit_it_17_vnu_189_in_2, msg_to_bit_it_17_vnu_190_in_0, msg_to_bit_it_17_vnu_190_in_1, msg_to_bit_it_17_vnu_190_in_2, msg_to_bit_it_17_vnu_191_in_0, msg_to_bit_it_17_vnu_191_in_1, msg_to_bit_it_17_vnu_191_in_2, msg_to_bit_it_17_vnu_192_in_0, msg_to_bit_it_17_vnu_192_in_1, msg_to_bit_it_17_vnu_192_in_2, msg_to_bit_it_17_vnu_193_in_0, msg_to_bit_it_17_vnu_193_in_1, msg_to_bit_it_17_vnu_193_in_2, msg_to_bit_it_17_vnu_194_in_0, msg_to_bit_it_17_vnu_194_in_1, msg_to_bit_it_17_vnu_194_in_2, msg_to_bit_it_17_vnu_195_in_0, msg_to_bit_it_17_vnu_195_in_1, msg_to_bit_it_17_vnu_195_in_2, msg_to_bit_it_17_vnu_196_in_0, msg_to_bit_it_17_vnu_196_in_1, msg_to_bit_it_17_vnu_196_in_2, msg_to_bit_it_17_vnu_197_in_0, msg_to_bit_it_17_vnu_197_in_1, msg_to_bit_it_17_vnu_197_in_2, msg_to_bit_it_18_vnu_0_in_0, msg_to_bit_it_18_vnu_0_in_1, msg_to_bit_it_18_vnu_0_in_2, msg_to_bit_it_18_vnu_1_in_0, msg_to_bit_it_18_vnu_1_in_1, msg_to_bit_it_18_vnu_1_in_2, msg_to_bit_it_18_vnu_2_in_0, msg_to_bit_it_18_vnu_2_in_1, msg_to_bit_it_18_vnu_2_in_2, msg_to_bit_it_18_vnu_3_in_0, msg_to_bit_it_18_vnu_3_in_1, msg_to_bit_it_18_vnu_3_in_2, msg_to_bit_it_18_vnu_4_in_0, msg_to_bit_it_18_vnu_4_in_1, msg_to_bit_it_18_vnu_4_in_2, msg_to_bit_it_18_vnu_5_in_0, msg_to_bit_it_18_vnu_5_in_1, msg_to_bit_it_18_vnu_5_in_2, msg_to_bit_it_18_vnu_6_in_0, msg_to_bit_it_18_vnu_6_in_1, msg_to_bit_it_18_vnu_6_in_2, msg_to_bit_it_18_vnu_7_in_0, msg_to_bit_it_18_vnu_7_in_1, msg_to_bit_it_18_vnu_7_in_2, msg_to_bit_it_18_vnu_8_in_0, msg_to_bit_it_18_vnu_8_in_1, msg_to_bit_it_18_vnu_8_in_2, msg_to_bit_it_18_vnu_9_in_0, msg_to_bit_it_18_vnu_9_in_1, msg_to_bit_it_18_vnu_9_in_2, msg_to_bit_it_18_vnu_10_in_0, msg_to_bit_it_18_vnu_10_in_1, msg_to_bit_it_18_vnu_10_in_2, msg_to_bit_it_18_vnu_11_in_0, msg_to_bit_it_18_vnu_11_in_1, msg_to_bit_it_18_vnu_11_in_2, msg_to_bit_it_18_vnu_12_in_0, msg_to_bit_it_18_vnu_12_in_1, msg_to_bit_it_18_vnu_12_in_2, msg_to_bit_it_18_vnu_13_in_0, msg_to_bit_it_18_vnu_13_in_1, msg_to_bit_it_18_vnu_13_in_2, msg_to_bit_it_18_vnu_14_in_0, msg_to_bit_it_18_vnu_14_in_1, msg_to_bit_it_18_vnu_14_in_2, msg_to_bit_it_18_vnu_15_in_0, msg_to_bit_it_18_vnu_15_in_1, msg_to_bit_it_18_vnu_15_in_2, msg_to_bit_it_18_vnu_16_in_0, msg_to_bit_it_18_vnu_16_in_1, msg_to_bit_it_18_vnu_16_in_2, msg_to_bit_it_18_vnu_17_in_0, msg_to_bit_it_18_vnu_17_in_1, msg_to_bit_it_18_vnu_17_in_2, msg_to_bit_it_18_vnu_18_in_0, msg_to_bit_it_18_vnu_18_in_1, msg_to_bit_it_18_vnu_18_in_2, msg_to_bit_it_18_vnu_19_in_0, msg_to_bit_it_18_vnu_19_in_1, msg_to_bit_it_18_vnu_19_in_2, msg_to_bit_it_18_vnu_20_in_0, msg_to_bit_it_18_vnu_20_in_1, msg_to_bit_it_18_vnu_20_in_2, msg_to_bit_it_18_vnu_21_in_0, msg_to_bit_it_18_vnu_21_in_1, msg_to_bit_it_18_vnu_21_in_2, msg_to_bit_it_18_vnu_22_in_0, msg_to_bit_it_18_vnu_22_in_1, msg_to_bit_it_18_vnu_22_in_2, msg_to_bit_it_18_vnu_23_in_0, msg_to_bit_it_18_vnu_23_in_1, msg_to_bit_it_18_vnu_23_in_2, msg_to_bit_it_18_vnu_24_in_0, msg_to_bit_it_18_vnu_24_in_1, msg_to_bit_it_18_vnu_24_in_2, msg_to_bit_it_18_vnu_25_in_0, msg_to_bit_it_18_vnu_25_in_1, msg_to_bit_it_18_vnu_25_in_2, msg_to_bit_it_18_vnu_26_in_0, msg_to_bit_it_18_vnu_26_in_1, msg_to_bit_it_18_vnu_26_in_2, msg_to_bit_it_18_vnu_27_in_0, msg_to_bit_it_18_vnu_27_in_1, msg_to_bit_it_18_vnu_27_in_2, msg_to_bit_it_18_vnu_28_in_0, msg_to_bit_it_18_vnu_28_in_1, msg_to_bit_it_18_vnu_28_in_2, msg_to_bit_it_18_vnu_29_in_0, msg_to_bit_it_18_vnu_29_in_1, msg_to_bit_it_18_vnu_29_in_2, msg_to_bit_it_18_vnu_30_in_0, msg_to_bit_it_18_vnu_30_in_1, msg_to_bit_it_18_vnu_30_in_2, msg_to_bit_it_18_vnu_31_in_0, msg_to_bit_it_18_vnu_31_in_1, msg_to_bit_it_18_vnu_31_in_2, msg_to_bit_it_18_vnu_32_in_0, msg_to_bit_it_18_vnu_32_in_1, msg_to_bit_it_18_vnu_32_in_2, msg_to_bit_it_18_vnu_33_in_0, msg_to_bit_it_18_vnu_33_in_1, msg_to_bit_it_18_vnu_33_in_2, msg_to_bit_it_18_vnu_34_in_0, msg_to_bit_it_18_vnu_34_in_1, msg_to_bit_it_18_vnu_34_in_2, msg_to_bit_it_18_vnu_35_in_0, msg_to_bit_it_18_vnu_35_in_1, msg_to_bit_it_18_vnu_35_in_2, msg_to_bit_it_18_vnu_36_in_0, msg_to_bit_it_18_vnu_36_in_1, msg_to_bit_it_18_vnu_36_in_2, msg_to_bit_it_18_vnu_37_in_0, msg_to_bit_it_18_vnu_37_in_1, msg_to_bit_it_18_vnu_37_in_2, msg_to_bit_it_18_vnu_38_in_0, msg_to_bit_it_18_vnu_38_in_1, msg_to_bit_it_18_vnu_38_in_2, msg_to_bit_it_18_vnu_39_in_0, msg_to_bit_it_18_vnu_39_in_1, msg_to_bit_it_18_vnu_39_in_2, msg_to_bit_it_18_vnu_40_in_0, msg_to_bit_it_18_vnu_40_in_1, msg_to_bit_it_18_vnu_40_in_2, msg_to_bit_it_18_vnu_41_in_0, msg_to_bit_it_18_vnu_41_in_1, msg_to_bit_it_18_vnu_41_in_2, msg_to_bit_it_18_vnu_42_in_0, msg_to_bit_it_18_vnu_42_in_1, msg_to_bit_it_18_vnu_42_in_2, msg_to_bit_it_18_vnu_43_in_0, msg_to_bit_it_18_vnu_43_in_1, msg_to_bit_it_18_vnu_43_in_2, msg_to_bit_it_18_vnu_44_in_0, msg_to_bit_it_18_vnu_44_in_1, msg_to_bit_it_18_vnu_44_in_2, msg_to_bit_it_18_vnu_45_in_0, msg_to_bit_it_18_vnu_45_in_1, msg_to_bit_it_18_vnu_45_in_2, msg_to_bit_it_18_vnu_46_in_0, msg_to_bit_it_18_vnu_46_in_1, msg_to_bit_it_18_vnu_46_in_2, msg_to_bit_it_18_vnu_47_in_0, msg_to_bit_it_18_vnu_47_in_1, msg_to_bit_it_18_vnu_47_in_2, msg_to_bit_it_18_vnu_48_in_0, msg_to_bit_it_18_vnu_48_in_1, msg_to_bit_it_18_vnu_48_in_2, msg_to_bit_it_18_vnu_49_in_0, msg_to_bit_it_18_vnu_49_in_1, msg_to_bit_it_18_vnu_49_in_2, msg_to_bit_it_18_vnu_50_in_0, msg_to_bit_it_18_vnu_50_in_1, msg_to_bit_it_18_vnu_50_in_2, msg_to_bit_it_18_vnu_51_in_0, msg_to_bit_it_18_vnu_51_in_1, msg_to_bit_it_18_vnu_51_in_2, msg_to_bit_it_18_vnu_52_in_0, msg_to_bit_it_18_vnu_52_in_1, msg_to_bit_it_18_vnu_52_in_2, msg_to_bit_it_18_vnu_53_in_0, msg_to_bit_it_18_vnu_53_in_1, msg_to_bit_it_18_vnu_53_in_2, msg_to_bit_it_18_vnu_54_in_0, msg_to_bit_it_18_vnu_54_in_1, msg_to_bit_it_18_vnu_54_in_2, msg_to_bit_it_18_vnu_55_in_0, msg_to_bit_it_18_vnu_55_in_1, msg_to_bit_it_18_vnu_55_in_2, msg_to_bit_it_18_vnu_56_in_0, msg_to_bit_it_18_vnu_56_in_1, msg_to_bit_it_18_vnu_56_in_2, msg_to_bit_it_18_vnu_57_in_0, msg_to_bit_it_18_vnu_57_in_1, msg_to_bit_it_18_vnu_57_in_2, msg_to_bit_it_18_vnu_58_in_0, msg_to_bit_it_18_vnu_58_in_1, msg_to_bit_it_18_vnu_58_in_2, msg_to_bit_it_18_vnu_59_in_0, msg_to_bit_it_18_vnu_59_in_1, msg_to_bit_it_18_vnu_59_in_2, msg_to_bit_it_18_vnu_60_in_0, msg_to_bit_it_18_vnu_60_in_1, msg_to_bit_it_18_vnu_60_in_2, msg_to_bit_it_18_vnu_61_in_0, msg_to_bit_it_18_vnu_61_in_1, msg_to_bit_it_18_vnu_61_in_2, msg_to_bit_it_18_vnu_62_in_0, msg_to_bit_it_18_vnu_62_in_1, msg_to_bit_it_18_vnu_62_in_2, msg_to_bit_it_18_vnu_63_in_0, msg_to_bit_it_18_vnu_63_in_1, msg_to_bit_it_18_vnu_63_in_2, msg_to_bit_it_18_vnu_64_in_0, msg_to_bit_it_18_vnu_64_in_1, msg_to_bit_it_18_vnu_64_in_2, msg_to_bit_it_18_vnu_65_in_0, msg_to_bit_it_18_vnu_65_in_1, msg_to_bit_it_18_vnu_65_in_2, msg_to_bit_it_18_vnu_66_in_0, msg_to_bit_it_18_vnu_66_in_1, msg_to_bit_it_18_vnu_66_in_2, msg_to_bit_it_18_vnu_67_in_0, msg_to_bit_it_18_vnu_67_in_1, msg_to_bit_it_18_vnu_67_in_2, msg_to_bit_it_18_vnu_68_in_0, msg_to_bit_it_18_vnu_68_in_1, msg_to_bit_it_18_vnu_68_in_2, msg_to_bit_it_18_vnu_69_in_0, msg_to_bit_it_18_vnu_69_in_1, msg_to_bit_it_18_vnu_69_in_2, msg_to_bit_it_18_vnu_70_in_0, msg_to_bit_it_18_vnu_70_in_1, msg_to_bit_it_18_vnu_70_in_2, msg_to_bit_it_18_vnu_71_in_0, msg_to_bit_it_18_vnu_71_in_1, msg_to_bit_it_18_vnu_71_in_2, msg_to_bit_it_18_vnu_72_in_0, msg_to_bit_it_18_vnu_72_in_1, msg_to_bit_it_18_vnu_72_in_2, msg_to_bit_it_18_vnu_73_in_0, msg_to_bit_it_18_vnu_73_in_1, msg_to_bit_it_18_vnu_73_in_2, msg_to_bit_it_18_vnu_74_in_0, msg_to_bit_it_18_vnu_74_in_1, msg_to_bit_it_18_vnu_74_in_2, msg_to_bit_it_18_vnu_75_in_0, msg_to_bit_it_18_vnu_75_in_1, msg_to_bit_it_18_vnu_75_in_2, msg_to_bit_it_18_vnu_76_in_0, msg_to_bit_it_18_vnu_76_in_1, msg_to_bit_it_18_vnu_76_in_2, msg_to_bit_it_18_vnu_77_in_0, msg_to_bit_it_18_vnu_77_in_1, msg_to_bit_it_18_vnu_77_in_2, msg_to_bit_it_18_vnu_78_in_0, msg_to_bit_it_18_vnu_78_in_1, msg_to_bit_it_18_vnu_78_in_2, msg_to_bit_it_18_vnu_79_in_0, msg_to_bit_it_18_vnu_79_in_1, msg_to_bit_it_18_vnu_79_in_2, msg_to_bit_it_18_vnu_80_in_0, msg_to_bit_it_18_vnu_80_in_1, msg_to_bit_it_18_vnu_80_in_2, msg_to_bit_it_18_vnu_81_in_0, msg_to_bit_it_18_vnu_81_in_1, msg_to_bit_it_18_vnu_81_in_2, msg_to_bit_it_18_vnu_82_in_0, msg_to_bit_it_18_vnu_82_in_1, msg_to_bit_it_18_vnu_82_in_2, msg_to_bit_it_18_vnu_83_in_0, msg_to_bit_it_18_vnu_83_in_1, msg_to_bit_it_18_vnu_83_in_2, msg_to_bit_it_18_vnu_84_in_0, msg_to_bit_it_18_vnu_84_in_1, msg_to_bit_it_18_vnu_84_in_2, msg_to_bit_it_18_vnu_85_in_0, msg_to_bit_it_18_vnu_85_in_1, msg_to_bit_it_18_vnu_85_in_2, msg_to_bit_it_18_vnu_86_in_0, msg_to_bit_it_18_vnu_86_in_1, msg_to_bit_it_18_vnu_86_in_2, msg_to_bit_it_18_vnu_87_in_0, msg_to_bit_it_18_vnu_87_in_1, msg_to_bit_it_18_vnu_87_in_2, msg_to_bit_it_18_vnu_88_in_0, msg_to_bit_it_18_vnu_88_in_1, msg_to_bit_it_18_vnu_88_in_2, msg_to_bit_it_18_vnu_89_in_0, msg_to_bit_it_18_vnu_89_in_1, msg_to_bit_it_18_vnu_89_in_2, msg_to_bit_it_18_vnu_90_in_0, msg_to_bit_it_18_vnu_90_in_1, msg_to_bit_it_18_vnu_90_in_2, msg_to_bit_it_18_vnu_91_in_0, msg_to_bit_it_18_vnu_91_in_1, msg_to_bit_it_18_vnu_91_in_2, msg_to_bit_it_18_vnu_92_in_0, msg_to_bit_it_18_vnu_92_in_1, msg_to_bit_it_18_vnu_92_in_2, msg_to_bit_it_18_vnu_93_in_0, msg_to_bit_it_18_vnu_93_in_1, msg_to_bit_it_18_vnu_93_in_2, msg_to_bit_it_18_vnu_94_in_0, msg_to_bit_it_18_vnu_94_in_1, msg_to_bit_it_18_vnu_94_in_2, msg_to_bit_it_18_vnu_95_in_0, msg_to_bit_it_18_vnu_95_in_1, msg_to_bit_it_18_vnu_95_in_2, msg_to_bit_it_18_vnu_96_in_0, msg_to_bit_it_18_vnu_96_in_1, msg_to_bit_it_18_vnu_96_in_2, msg_to_bit_it_18_vnu_97_in_0, msg_to_bit_it_18_vnu_97_in_1, msg_to_bit_it_18_vnu_97_in_2, msg_to_bit_it_18_vnu_98_in_0, msg_to_bit_it_18_vnu_98_in_1, msg_to_bit_it_18_vnu_98_in_2, msg_to_bit_it_18_vnu_99_in_0, msg_to_bit_it_18_vnu_99_in_1, msg_to_bit_it_18_vnu_99_in_2, msg_to_bit_it_18_vnu_100_in_0, msg_to_bit_it_18_vnu_100_in_1, msg_to_bit_it_18_vnu_100_in_2, msg_to_bit_it_18_vnu_101_in_0, msg_to_bit_it_18_vnu_101_in_1, msg_to_bit_it_18_vnu_101_in_2, msg_to_bit_it_18_vnu_102_in_0, msg_to_bit_it_18_vnu_102_in_1, msg_to_bit_it_18_vnu_102_in_2, msg_to_bit_it_18_vnu_103_in_0, msg_to_bit_it_18_vnu_103_in_1, msg_to_bit_it_18_vnu_103_in_2, msg_to_bit_it_18_vnu_104_in_0, msg_to_bit_it_18_vnu_104_in_1, msg_to_bit_it_18_vnu_104_in_2, msg_to_bit_it_18_vnu_105_in_0, msg_to_bit_it_18_vnu_105_in_1, msg_to_bit_it_18_vnu_105_in_2, msg_to_bit_it_18_vnu_106_in_0, msg_to_bit_it_18_vnu_106_in_1, msg_to_bit_it_18_vnu_106_in_2, msg_to_bit_it_18_vnu_107_in_0, msg_to_bit_it_18_vnu_107_in_1, msg_to_bit_it_18_vnu_107_in_2, msg_to_bit_it_18_vnu_108_in_0, msg_to_bit_it_18_vnu_108_in_1, msg_to_bit_it_18_vnu_108_in_2, msg_to_bit_it_18_vnu_109_in_0, msg_to_bit_it_18_vnu_109_in_1, msg_to_bit_it_18_vnu_109_in_2, msg_to_bit_it_18_vnu_110_in_0, msg_to_bit_it_18_vnu_110_in_1, msg_to_bit_it_18_vnu_110_in_2, msg_to_bit_it_18_vnu_111_in_0, msg_to_bit_it_18_vnu_111_in_1, msg_to_bit_it_18_vnu_111_in_2, msg_to_bit_it_18_vnu_112_in_0, msg_to_bit_it_18_vnu_112_in_1, msg_to_bit_it_18_vnu_112_in_2, msg_to_bit_it_18_vnu_113_in_0, msg_to_bit_it_18_vnu_113_in_1, msg_to_bit_it_18_vnu_113_in_2, msg_to_bit_it_18_vnu_114_in_0, msg_to_bit_it_18_vnu_114_in_1, msg_to_bit_it_18_vnu_114_in_2, msg_to_bit_it_18_vnu_115_in_0, msg_to_bit_it_18_vnu_115_in_1, msg_to_bit_it_18_vnu_115_in_2, msg_to_bit_it_18_vnu_116_in_0, msg_to_bit_it_18_vnu_116_in_1, msg_to_bit_it_18_vnu_116_in_2, msg_to_bit_it_18_vnu_117_in_0, msg_to_bit_it_18_vnu_117_in_1, msg_to_bit_it_18_vnu_117_in_2, msg_to_bit_it_18_vnu_118_in_0, msg_to_bit_it_18_vnu_118_in_1, msg_to_bit_it_18_vnu_118_in_2, msg_to_bit_it_18_vnu_119_in_0, msg_to_bit_it_18_vnu_119_in_1, msg_to_bit_it_18_vnu_119_in_2, msg_to_bit_it_18_vnu_120_in_0, msg_to_bit_it_18_vnu_120_in_1, msg_to_bit_it_18_vnu_120_in_2, msg_to_bit_it_18_vnu_121_in_0, msg_to_bit_it_18_vnu_121_in_1, msg_to_bit_it_18_vnu_121_in_2, msg_to_bit_it_18_vnu_122_in_0, msg_to_bit_it_18_vnu_122_in_1, msg_to_bit_it_18_vnu_122_in_2, msg_to_bit_it_18_vnu_123_in_0, msg_to_bit_it_18_vnu_123_in_1, msg_to_bit_it_18_vnu_123_in_2, msg_to_bit_it_18_vnu_124_in_0, msg_to_bit_it_18_vnu_124_in_1, msg_to_bit_it_18_vnu_124_in_2, msg_to_bit_it_18_vnu_125_in_0, msg_to_bit_it_18_vnu_125_in_1, msg_to_bit_it_18_vnu_125_in_2, msg_to_bit_it_18_vnu_126_in_0, msg_to_bit_it_18_vnu_126_in_1, msg_to_bit_it_18_vnu_126_in_2, msg_to_bit_it_18_vnu_127_in_0, msg_to_bit_it_18_vnu_127_in_1, msg_to_bit_it_18_vnu_127_in_2, msg_to_bit_it_18_vnu_128_in_0, msg_to_bit_it_18_vnu_128_in_1, msg_to_bit_it_18_vnu_128_in_2, msg_to_bit_it_18_vnu_129_in_0, msg_to_bit_it_18_vnu_129_in_1, msg_to_bit_it_18_vnu_129_in_2, msg_to_bit_it_18_vnu_130_in_0, msg_to_bit_it_18_vnu_130_in_1, msg_to_bit_it_18_vnu_130_in_2, msg_to_bit_it_18_vnu_131_in_0, msg_to_bit_it_18_vnu_131_in_1, msg_to_bit_it_18_vnu_131_in_2, msg_to_bit_it_18_vnu_132_in_0, msg_to_bit_it_18_vnu_132_in_1, msg_to_bit_it_18_vnu_132_in_2, msg_to_bit_it_18_vnu_133_in_0, msg_to_bit_it_18_vnu_133_in_1, msg_to_bit_it_18_vnu_133_in_2, msg_to_bit_it_18_vnu_134_in_0, msg_to_bit_it_18_vnu_134_in_1, msg_to_bit_it_18_vnu_134_in_2, msg_to_bit_it_18_vnu_135_in_0, msg_to_bit_it_18_vnu_135_in_1, msg_to_bit_it_18_vnu_135_in_2, msg_to_bit_it_18_vnu_136_in_0, msg_to_bit_it_18_vnu_136_in_1, msg_to_bit_it_18_vnu_136_in_2, msg_to_bit_it_18_vnu_137_in_0, msg_to_bit_it_18_vnu_137_in_1, msg_to_bit_it_18_vnu_137_in_2, msg_to_bit_it_18_vnu_138_in_0, msg_to_bit_it_18_vnu_138_in_1, msg_to_bit_it_18_vnu_138_in_2, msg_to_bit_it_18_vnu_139_in_0, msg_to_bit_it_18_vnu_139_in_1, msg_to_bit_it_18_vnu_139_in_2, msg_to_bit_it_18_vnu_140_in_0, msg_to_bit_it_18_vnu_140_in_1, msg_to_bit_it_18_vnu_140_in_2, msg_to_bit_it_18_vnu_141_in_0, msg_to_bit_it_18_vnu_141_in_1, msg_to_bit_it_18_vnu_141_in_2, msg_to_bit_it_18_vnu_142_in_0, msg_to_bit_it_18_vnu_142_in_1, msg_to_bit_it_18_vnu_142_in_2, msg_to_bit_it_18_vnu_143_in_0, msg_to_bit_it_18_vnu_143_in_1, msg_to_bit_it_18_vnu_143_in_2, msg_to_bit_it_18_vnu_144_in_0, msg_to_bit_it_18_vnu_144_in_1, msg_to_bit_it_18_vnu_144_in_2, msg_to_bit_it_18_vnu_145_in_0, msg_to_bit_it_18_vnu_145_in_1, msg_to_bit_it_18_vnu_145_in_2, msg_to_bit_it_18_vnu_146_in_0, msg_to_bit_it_18_vnu_146_in_1, msg_to_bit_it_18_vnu_146_in_2, msg_to_bit_it_18_vnu_147_in_0, msg_to_bit_it_18_vnu_147_in_1, msg_to_bit_it_18_vnu_147_in_2, msg_to_bit_it_18_vnu_148_in_0, msg_to_bit_it_18_vnu_148_in_1, msg_to_bit_it_18_vnu_148_in_2, msg_to_bit_it_18_vnu_149_in_0, msg_to_bit_it_18_vnu_149_in_1, msg_to_bit_it_18_vnu_149_in_2, msg_to_bit_it_18_vnu_150_in_0, msg_to_bit_it_18_vnu_150_in_1, msg_to_bit_it_18_vnu_150_in_2, msg_to_bit_it_18_vnu_151_in_0, msg_to_bit_it_18_vnu_151_in_1, msg_to_bit_it_18_vnu_151_in_2, msg_to_bit_it_18_vnu_152_in_0, msg_to_bit_it_18_vnu_152_in_1, msg_to_bit_it_18_vnu_152_in_2, msg_to_bit_it_18_vnu_153_in_0, msg_to_bit_it_18_vnu_153_in_1, msg_to_bit_it_18_vnu_153_in_2, msg_to_bit_it_18_vnu_154_in_0, msg_to_bit_it_18_vnu_154_in_1, msg_to_bit_it_18_vnu_154_in_2, msg_to_bit_it_18_vnu_155_in_0, msg_to_bit_it_18_vnu_155_in_1, msg_to_bit_it_18_vnu_155_in_2, msg_to_bit_it_18_vnu_156_in_0, msg_to_bit_it_18_vnu_156_in_1, msg_to_bit_it_18_vnu_156_in_2, msg_to_bit_it_18_vnu_157_in_0, msg_to_bit_it_18_vnu_157_in_1, msg_to_bit_it_18_vnu_157_in_2, msg_to_bit_it_18_vnu_158_in_0, msg_to_bit_it_18_vnu_158_in_1, msg_to_bit_it_18_vnu_158_in_2, msg_to_bit_it_18_vnu_159_in_0, msg_to_bit_it_18_vnu_159_in_1, msg_to_bit_it_18_vnu_159_in_2, msg_to_bit_it_18_vnu_160_in_0, msg_to_bit_it_18_vnu_160_in_1, msg_to_bit_it_18_vnu_160_in_2, msg_to_bit_it_18_vnu_161_in_0, msg_to_bit_it_18_vnu_161_in_1, msg_to_bit_it_18_vnu_161_in_2, msg_to_bit_it_18_vnu_162_in_0, msg_to_bit_it_18_vnu_162_in_1, msg_to_bit_it_18_vnu_162_in_2, msg_to_bit_it_18_vnu_163_in_0, msg_to_bit_it_18_vnu_163_in_1, msg_to_bit_it_18_vnu_163_in_2, msg_to_bit_it_18_vnu_164_in_0, msg_to_bit_it_18_vnu_164_in_1, msg_to_bit_it_18_vnu_164_in_2, msg_to_bit_it_18_vnu_165_in_0, msg_to_bit_it_18_vnu_165_in_1, msg_to_bit_it_18_vnu_165_in_2, msg_to_bit_it_18_vnu_166_in_0, msg_to_bit_it_18_vnu_166_in_1, msg_to_bit_it_18_vnu_166_in_2, msg_to_bit_it_18_vnu_167_in_0, msg_to_bit_it_18_vnu_167_in_1, msg_to_bit_it_18_vnu_167_in_2, msg_to_bit_it_18_vnu_168_in_0, msg_to_bit_it_18_vnu_168_in_1, msg_to_bit_it_18_vnu_168_in_2, msg_to_bit_it_18_vnu_169_in_0, msg_to_bit_it_18_vnu_169_in_1, msg_to_bit_it_18_vnu_169_in_2, msg_to_bit_it_18_vnu_170_in_0, msg_to_bit_it_18_vnu_170_in_1, msg_to_bit_it_18_vnu_170_in_2, msg_to_bit_it_18_vnu_171_in_0, msg_to_bit_it_18_vnu_171_in_1, msg_to_bit_it_18_vnu_171_in_2, msg_to_bit_it_18_vnu_172_in_0, msg_to_bit_it_18_vnu_172_in_1, msg_to_bit_it_18_vnu_172_in_2, msg_to_bit_it_18_vnu_173_in_0, msg_to_bit_it_18_vnu_173_in_1, msg_to_bit_it_18_vnu_173_in_2, msg_to_bit_it_18_vnu_174_in_0, msg_to_bit_it_18_vnu_174_in_1, msg_to_bit_it_18_vnu_174_in_2, msg_to_bit_it_18_vnu_175_in_0, msg_to_bit_it_18_vnu_175_in_1, msg_to_bit_it_18_vnu_175_in_2, msg_to_bit_it_18_vnu_176_in_0, msg_to_bit_it_18_vnu_176_in_1, msg_to_bit_it_18_vnu_176_in_2, msg_to_bit_it_18_vnu_177_in_0, msg_to_bit_it_18_vnu_177_in_1, msg_to_bit_it_18_vnu_177_in_2, msg_to_bit_it_18_vnu_178_in_0, msg_to_bit_it_18_vnu_178_in_1, msg_to_bit_it_18_vnu_178_in_2, msg_to_bit_it_18_vnu_179_in_0, msg_to_bit_it_18_vnu_179_in_1, msg_to_bit_it_18_vnu_179_in_2, msg_to_bit_it_18_vnu_180_in_0, msg_to_bit_it_18_vnu_180_in_1, msg_to_bit_it_18_vnu_180_in_2, msg_to_bit_it_18_vnu_181_in_0, msg_to_bit_it_18_vnu_181_in_1, msg_to_bit_it_18_vnu_181_in_2, msg_to_bit_it_18_vnu_182_in_0, msg_to_bit_it_18_vnu_182_in_1, msg_to_bit_it_18_vnu_182_in_2, msg_to_bit_it_18_vnu_183_in_0, msg_to_bit_it_18_vnu_183_in_1, msg_to_bit_it_18_vnu_183_in_2, msg_to_bit_it_18_vnu_184_in_0, msg_to_bit_it_18_vnu_184_in_1, msg_to_bit_it_18_vnu_184_in_2, msg_to_bit_it_18_vnu_185_in_0, msg_to_bit_it_18_vnu_185_in_1, msg_to_bit_it_18_vnu_185_in_2, msg_to_bit_it_18_vnu_186_in_0, msg_to_bit_it_18_vnu_186_in_1, msg_to_bit_it_18_vnu_186_in_2, msg_to_bit_it_18_vnu_187_in_0, msg_to_bit_it_18_vnu_187_in_1, msg_to_bit_it_18_vnu_187_in_2, msg_to_bit_it_18_vnu_188_in_0, msg_to_bit_it_18_vnu_188_in_1, msg_to_bit_it_18_vnu_188_in_2, msg_to_bit_it_18_vnu_189_in_0, msg_to_bit_it_18_vnu_189_in_1, msg_to_bit_it_18_vnu_189_in_2, msg_to_bit_it_18_vnu_190_in_0, msg_to_bit_it_18_vnu_190_in_1, msg_to_bit_it_18_vnu_190_in_2, msg_to_bit_it_18_vnu_191_in_0, msg_to_bit_it_18_vnu_191_in_1, msg_to_bit_it_18_vnu_191_in_2, msg_to_bit_it_18_vnu_192_in_0, msg_to_bit_it_18_vnu_192_in_1, msg_to_bit_it_18_vnu_192_in_2, msg_to_bit_it_18_vnu_193_in_0, msg_to_bit_it_18_vnu_193_in_1, msg_to_bit_it_18_vnu_193_in_2, msg_to_bit_it_18_vnu_194_in_0, msg_to_bit_it_18_vnu_194_in_1, msg_to_bit_it_18_vnu_194_in_2, msg_to_bit_it_18_vnu_195_in_0, msg_to_bit_it_18_vnu_195_in_1, msg_to_bit_it_18_vnu_195_in_2, msg_to_bit_it_18_vnu_196_in_0, msg_to_bit_it_18_vnu_196_in_1, msg_to_bit_it_18_vnu_196_in_2, msg_to_bit_it_18_vnu_197_in_0, msg_to_bit_it_18_vnu_197_in_1, msg_to_bit_it_18_vnu_197_in_2, msg_to_bit_it_19_vnu_0_in_0, msg_to_bit_it_19_vnu_0_in_1, msg_to_bit_it_19_vnu_0_in_2, msg_to_bit_it_19_vnu_1_in_0, msg_to_bit_it_19_vnu_1_in_1, msg_to_bit_it_19_vnu_1_in_2, msg_to_bit_it_19_vnu_2_in_0, msg_to_bit_it_19_vnu_2_in_1, msg_to_bit_it_19_vnu_2_in_2, msg_to_bit_it_19_vnu_3_in_0, msg_to_bit_it_19_vnu_3_in_1, msg_to_bit_it_19_vnu_3_in_2, msg_to_bit_it_19_vnu_4_in_0, msg_to_bit_it_19_vnu_4_in_1, msg_to_bit_it_19_vnu_4_in_2, msg_to_bit_it_19_vnu_5_in_0, msg_to_bit_it_19_vnu_5_in_1, msg_to_bit_it_19_vnu_5_in_2, msg_to_bit_it_19_vnu_6_in_0, msg_to_bit_it_19_vnu_6_in_1, msg_to_bit_it_19_vnu_6_in_2, msg_to_bit_it_19_vnu_7_in_0, msg_to_bit_it_19_vnu_7_in_1, msg_to_bit_it_19_vnu_7_in_2, msg_to_bit_it_19_vnu_8_in_0, msg_to_bit_it_19_vnu_8_in_1, msg_to_bit_it_19_vnu_8_in_2, msg_to_bit_it_19_vnu_9_in_0, msg_to_bit_it_19_vnu_9_in_1, msg_to_bit_it_19_vnu_9_in_2, msg_to_bit_it_19_vnu_10_in_0, msg_to_bit_it_19_vnu_10_in_1, msg_to_bit_it_19_vnu_10_in_2, msg_to_bit_it_19_vnu_11_in_0, msg_to_bit_it_19_vnu_11_in_1, msg_to_bit_it_19_vnu_11_in_2, msg_to_bit_it_19_vnu_12_in_0, msg_to_bit_it_19_vnu_12_in_1, msg_to_bit_it_19_vnu_12_in_2, msg_to_bit_it_19_vnu_13_in_0, msg_to_bit_it_19_vnu_13_in_1, msg_to_bit_it_19_vnu_13_in_2, msg_to_bit_it_19_vnu_14_in_0, msg_to_bit_it_19_vnu_14_in_1, msg_to_bit_it_19_vnu_14_in_2, msg_to_bit_it_19_vnu_15_in_0, msg_to_bit_it_19_vnu_15_in_1, msg_to_bit_it_19_vnu_15_in_2, msg_to_bit_it_19_vnu_16_in_0, msg_to_bit_it_19_vnu_16_in_1, msg_to_bit_it_19_vnu_16_in_2, msg_to_bit_it_19_vnu_17_in_0, msg_to_bit_it_19_vnu_17_in_1, msg_to_bit_it_19_vnu_17_in_2, msg_to_bit_it_19_vnu_18_in_0, msg_to_bit_it_19_vnu_18_in_1, msg_to_bit_it_19_vnu_18_in_2, msg_to_bit_it_19_vnu_19_in_0, msg_to_bit_it_19_vnu_19_in_1, msg_to_bit_it_19_vnu_19_in_2, msg_to_bit_it_19_vnu_20_in_0, msg_to_bit_it_19_vnu_20_in_1, msg_to_bit_it_19_vnu_20_in_2, msg_to_bit_it_19_vnu_21_in_0, msg_to_bit_it_19_vnu_21_in_1, msg_to_bit_it_19_vnu_21_in_2, msg_to_bit_it_19_vnu_22_in_0, msg_to_bit_it_19_vnu_22_in_1, msg_to_bit_it_19_vnu_22_in_2, msg_to_bit_it_19_vnu_23_in_0, msg_to_bit_it_19_vnu_23_in_1, msg_to_bit_it_19_vnu_23_in_2, msg_to_bit_it_19_vnu_24_in_0, msg_to_bit_it_19_vnu_24_in_1, msg_to_bit_it_19_vnu_24_in_2, msg_to_bit_it_19_vnu_25_in_0, msg_to_bit_it_19_vnu_25_in_1, msg_to_bit_it_19_vnu_25_in_2, msg_to_bit_it_19_vnu_26_in_0, msg_to_bit_it_19_vnu_26_in_1, msg_to_bit_it_19_vnu_26_in_2, msg_to_bit_it_19_vnu_27_in_0, msg_to_bit_it_19_vnu_27_in_1, msg_to_bit_it_19_vnu_27_in_2, msg_to_bit_it_19_vnu_28_in_0, msg_to_bit_it_19_vnu_28_in_1, msg_to_bit_it_19_vnu_28_in_2, msg_to_bit_it_19_vnu_29_in_0, msg_to_bit_it_19_vnu_29_in_1, msg_to_bit_it_19_vnu_29_in_2, msg_to_bit_it_19_vnu_30_in_0, msg_to_bit_it_19_vnu_30_in_1, msg_to_bit_it_19_vnu_30_in_2, msg_to_bit_it_19_vnu_31_in_0, msg_to_bit_it_19_vnu_31_in_1, msg_to_bit_it_19_vnu_31_in_2, msg_to_bit_it_19_vnu_32_in_0, msg_to_bit_it_19_vnu_32_in_1, msg_to_bit_it_19_vnu_32_in_2, msg_to_bit_it_19_vnu_33_in_0, msg_to_bit_it_19_vnu_33_in_1, msg_to_bit_it_19_vnu_33_in_2, msg_to_bit_it_19_vnu_34_in_0, msg_to_bit_it_19_vnu_34_in_1, msg_to_bit_it_19_vnu_34_in_2, msg_to_bit_it_19_vnu_35_in_0, msg_to_bit_it_19_vnu_35_in_1, msg_to_bit_it_19_vnu_35_in_2, msg_to_bit_it_19_vnu_36_in_0, msg_to_bit_it_19_vnu_36_in_1, msg_to_bit_it_19_vnu_36_in_2, msg_to_bit_it_19_vnu_37_in_0, msg_to_bit_it_19_vnu_37_in_1, msg_to_bit_it_19_vnu_37_in_2, msg_to_bit_it_19_vnu_38_in_0, msg_to_bit_it_19_vnu_38_in_1, msg_to_bit_it_19_vnu_38_in_2, msg_to_bit_it_19_vnu_39_in_0, msg_to_bit_it_19_vnu_39_in_1, msg_to_bit_it_19_vnu_39_in_2, msg_to_bit_it_19_vnu_40_in_0, msg_to_bit_it_19_vnu_40_in_1, msg_to_bit_it_19_vnu_40_in_2, msg_to_bit_it_19_vnu_41_in_0, msg_to_bit_it_19_vnu_41_in_1, msg_to_bit_it_19_vnu_41_in_2, msg_to_bit_it_19_vnu_42_in_0, msg_to_bit_it_19_vnu_42_in_1, msg_to_bit_it_19_vnu_42_in_2, msg_to_bit_it_19_vnu_43_in_0, msg_to_bit_it_19_vnu_43_in_1, msg_to_bit_it_19_vnu_43_in_2, msg_to_bit_it_19_vnu_44_in_0, msg_to_bit_it_19_vnu_44_in_1, msg_to_bit_it_19_vnu_44_in_2, msg_to_bit_it_19_vnu_45_in_0, msg_to_bit_it_19_vnu_45_in_1, msg_to_bit_it_19_vnu_45_in_2, msg_to_bit_it_19_vnu_46_in_0, msg_to_bit_it_19_vnu_46_in_1, msg_to_bit_it_19_vnu_46_in_2, msg_to_bit_it_19_vnu_47_in_0, msg_to_bit_it_19_vnu_47_in_1, msg_to_bit_it_19_vnu_47_in_2, msg_to_bit_it_19_vnu_48_in_0, msg_to_bit_it_19_vnu_48_in_1, msg_to_bit_it_19_vnu_48_in_2, msg_to_bit_it_19_vnu_49_in_0, msg_to_bit_it_19_vnu_49_in_1, msg_to_bit_it_19_vnu_49_in_2, msg_to_bit_it_19_vnu_50_in_0, msg_to_bit_it_19_vnu_50_in_1, msg_to_bit_it_19_vnu_50_in_2, msg_to_bit_it_19_vnu_51_in_0, msg_to_bit_it_19_vnu_51_in_1, msg_to_bit_it_19_vnu_51_in_2, msg_to_bit_it_19_vnu_52_in_0, msg_to_bit_it_19_vnu_52_in_1, msg_to_bit_it_19_vnu_52_in_2, msg_to_bit_it_19_vnu_53_in_0, msg_to_bit_it_19_vnu_53_in_1, msg_to_bit_it_19_vnu_53_in_2, msg_to_bit_it_19_vnu_54_in_0, msg_to_bit_it_19_vnu_54_in_1, msg_to_bit_it_19_vnu_54_in_2, msg_to_bit_it_19_vnu_55_in_0, msg_to_bit_it_19_vnu_55_in_1, msg_to_bit_it_19_vnu_55_in_2, msg_to_bit_it_19_vnu_56_in_0, msg_to_bit_it_19_vnu_56_in_1, msg_to_bit_it_19_vnu_56_in_2, msg_to_bit_it_19_vnu_57_in_0, msg_to_bit_it_19_vnu_57_in_1, msg_to_bit_it_19_vnu_57_in_2, msg_to_bit_it_19_vnu_58_in_0, msg_to_bit_it_19_vnu_58_in_1, msg_to_bit_it_19_vnu_58_in_2, msg_to_bit_it_19_vnu_59_in_0, msg_to_bit_it_19_vnu_59_in_1, msg_to_bit_it_19_vnu_59_in_2, msg_to_bit_it_19_vnu_60_in_0, msg_to_bit_it_19_vnu_60_in_1, msg_to_bit_it_19_vnu_60_in_2, msg_to_bit_it_19_vnu_61_in_0, msg_to_bit_it_19_vnu_61_in_1, msg_to_bit_it_19_vnu_61_in_2, msg_to_bit_it_19_vnu_62_in_0, msg_to_bit_it_19_vnu_62_in_1, msg_to_bit_it_19_vnu_62_in_2, msg_to_bit_it_19_vnu_63_in_0, msg_to_bit_it_19_vnu_63_in_1, msg_to_bit_it_19_vnu_63_in_2, msg_to_bit_it_19_vnu_64_in_0, msg_to_bit_it_19_vnu_64_in_1, msg_to_bit_it_19_vnu_64_in_2, msg_to_bit_it_19_vnu_65_in_0, msg_to_bit_it_19_vnu_65_in_1, msg_to_bit_it_19_vnu_65_in_2, msg_to_bit_it_19_vnu_66_in_0, msg_to_bit_it_19_vnu_66_in_1, msg_to_bit_it_19_vnu_66_in_2, msg_to_bit_it_19_vnu_67_in_0, msg_to_bit_it_19_vnu_67_in_1, msg_to_bit_it_19_vnu_67_in_2, msg_to_bit_it_19_vnu_68_in_0, msg_to_bit_it_19_vnu_68_in_1, msg_to_bit_it_19_vnu_68_in_2, msg_to_bit_it_19_vnu_69_in_0, msg_to_bit_it_19_vnu_69_in_1, msg_to_bit_it_19_vnu_69_in_2, msg_to_bit_it_19_vnu_70_in_0, msg_to_bit_it_19_vnu_70_in_1, msg_to_bit_it_19_vnu_70_in_2, msg_to_bit_it_19_vnu_71_in_0, msg_to_bit_it_19_vnu_71_in_1, msg_to_bit_it_19_vnu_71_in_2, msg_to_bit_it_19_vnu_72_in_0, msg_to_bit_it_19_vnu_72_in_1, msg_to_bit_it_19_vnu_72_in_2, msg_to_bit_it_19_vnu_73_in_0, msg_to_bit_it_19_vnu_73_in_1, msg_to_bit_it_19_vnu_73_in_2, msg_to_bit_it_19_vnu_74_in_0, msg_to_bit_it_19_vnu_74_in_1, msg_to_bit_it_19_vnu_74_in_2, msg_to_bit_it_19_vnu_75_in_0, msg_to_bit_it_19_vnu_75_in_1, msg_to_bit_it_19_vnu_75_in_2, msg_to_bit_it_19_vnu_76_in_0, msg_to_bit_it_19_vnu_76_in_1, msg_to_bit_it_19_vnu_76_in_2, msg_to_bit_it_19_vnu_77_in_0, msg_to_bit_it_19_vnu_77_in_1, msg_to_bit_it_19_vnu_77_in_2, msg_to_bit_it_19_vnu_78_in_0, msg_to_bit_it_19_vnu_78_in_1, msg_to_bit_it_19_vnu_78_in_2, msg_to_bit_it_19_vnu_79_in_0, msg_to_bit_it_19_vnu_79_in_1, msg_to_bit_it_19_vnu_79_in_2, msg_to_bit_it_19_vnu_80_in_0, msg_to_bit_it_19_vnu_80_in_1, msg_to_bit_it_19_vnu_80_in_2, msg_to_bit_it_19_vnu_81_in_0, msg_to_bit_it_19_vnu_81_in_1, msg_to_bit_it_19_vnu_81_in_2, msg_to_bit_it_19_vnu_82_in_0, msg_to_bit_it_19_vnu_82_in_1, msg_to_bit_it_19_vnu_82_in_2, msg_to_bit_it_19_vnu_83_in_0, msg_to_bit_it_19_vnu_83_in_1, msg_to_bit_it_19_vnu_83_in_2, msg_to_bit_it_19_vnu_84_in_0, msg_to_bit_it_19_vnu_84_in_1, msg_to_bit_it_19_vnu_84_in_2, msg_to_bit_it_19_vnu_85_in_0, msg_to_bit_it_19_vnu_85_in_1, msg_to_bit_it_19_vnu_85_in_2, msg_to_bit_it_19_vnu_86_in_0, msg_to_bit_it_19_vnu_86_in_1, msg_to_bit_it_19_vnu_86_in_2, msg_to_bit_it_19_vnu_87_in_0, msg_to_bit_it_19_vnu_87_in_1, msg_to_bit_it_19_vnu_87_in_2, msg_to_bit_it_19_vnu_88_in_0, msg_to_bit_it_19_vnu_88_in_1, msg_to_bit_it_19_vnu_88_in_2, msg_to_bit_it_19_vnu_89_in_0, msg_to_bit_it_19_vnu_89_in_1, msg_to_bit_it_19_vnu_89_in_2, msg_to_bit_it_19_vnu_90_in_0, msg_to_bit_it_19_vnu_90_in_1, msg_to_bit_it_19_vnu_90_in_2, msg_to_bit_it_19_vnu_91_in_0, msg_to_bit_it_19_vnu_91_in_1, msg_to_bit_it_19_vnu_91_in_2, msg_to_bit_it_19_vnu_92_in_0, msg_to_bit_it_19_vnu_92_in_1, msg_to_bit_it_19_vnu_92_in_2, msg_to_bit_it_19_vnu_93_in_0, msg_to_bit_it_19_vnu_93_in_1, msg_to_bit_it_19_vnu_93_in_2, msg_to_bit_it_19_vnu_94_in_0, msg_to_bit_it_19_vnu_94_in_1, msg_to_bit_it_19_vnu_94_in_2, msg_to_bit_it_19_vnu_95_in_0, msg_to_bit_it_19_vnu_95_in_1, msg_to_bit_it_19_vnu_95_in_2, msg_to_bit_it_19_vnu_96_in_0, msg_to_bit_it_19_vnu_96_in_1, msg_to_bit_it_19_vnu_96_in_2, msg_to_bit_it_19_vnu_97_in_0, msg_to_bit_it_19_vnu_97_in_1, msg_to_bit_it_19_vnu_97_in_2, msg_to_bit_it_19_vnu_98_in_0, msg_to_bit_it_19_vnu_98_in_1, msg_to_bit_it_19_vnu_98_in_2, msg_to_bit_it_19_vnu_99_in_0, msg_to_bit_it_19_vnu_99_in_1, msg_to_bit_it_19_vnu_99_in_2, msg_to_bit_it_19_vnu_100_in_0, msg_to_bit_it_19_vnu_100_in_1, msg_to_bit_it_19_vnu_100_in_2, msg_to_bit_it_19_vnu_101_in_0, msg_to_bit_it_19_vnu_101_in_1, msg_to_bit_it_19_vnu_101_in_2, msg_to_bit_it_19_vnu_102_in_0, msg_to_bit_it_19_vnu_102_in_1, msg_to_bit_it_19_vnu_102_in_2, msg_to_bit_it_19_vnu_103_in_0, msg_to_bit_it_19_vnu_103_in_1, msg_to_bit_it_19_vnu_103_in_2, msg_to_bit_it_19_vnu_104_in_0, msg_to_bit_it_19_vnu_104_in_1, msg_to_bit_it_19_vnu_104_in_2, msg_to_bit_it_19_vnu_105_in_0, msg_to_bit_it_19_vnu_105_in_1, msg_to_bit_it_19_vnu_105_in_2, msg_to_bit_it_19_vnu_106_in_0, msg_to_bit_it_19_vnu_106_in_1, msg_to_bit_it_19_vnu_106_in_2, msg_to_bit_it_19_vnu_107_in_0, msg_to_bit_it_19_vnu_107_in_1, msg_to_bit_it_19_vnu_107_in_2, msg_to_bit_it_19_vnu_108_in_0, msg_to_bit_it_19_vnu_108_in_1, msg_to_bit_it_19_vnu_108_in_2, msg_to_bit_it_19_vnu_109_in_0, msg_to_bit_it_19_vnu_109_in_1, msg_to_bit_it_19_vnu_109_in_2, msg_to_bit_it_19_vnu_110_in_0, msg_to_bit_it_19_vnu_110_in_1, msg_to_bit_it_19_vnu_110_in_2, msg_to_bit_it_19_vnu_111_in_0, msg_to_bit_it_19_vnu_111_in_1, msg_to_bit_it_19_vnu_111_in_2, msg_to_bit_it_19_vnu_112_in_0, msg_to_bit_it_19_vnu_112_in_1, msg_to_bit_it_19_vnu_112_in_2, msg_to_bit_it_19_vnu_113_in_0, msg_to_bit_it_19_vnu_113_in_1, msg_to_bit_it_19_vnu_113_in_2, msg_to_bit_it_19_vnu_114_in_0, msg_to_bit_it_19_vnu_114_in_1, msg_to_bit_it_19_vnu_114_in_2, msg_to_bit_it_19_vnu_115_in_0, msg_to_bit_it_19_vnu_115_in_1, msg_to_bit_it_19_vnu_115_in_2, msg_to_bit_it_19_vnu_116_in_0, msg_to_bit_it_19_vnu_116_in_1, msg_to_bit_it_19_vnu_116_in_2, msg_to_bit_it_19_vnu_117_in_0, msg_to_bit_it_19_vnu_117_in_1, msg_to_bit_it_19_vnu_117_in_2, msg_to_bit_it_19_vnu_118_in_0, msg_to_bit_it_19_vnu_118_in_1, msg_to_bit_it_19_vnu_118_in_2, msg_to_bit_it_19_vnu_119_in_0, msg_to_bit_it_19_vnu_119_in_1, msg_to_bit_it_19_vnu_119_in_2, msg_to_bit_it_19_vnu_120_in_0, msg_to_bit_it_19_vnu_120_in_1, msg_to_bit_it_19_vnu_120_in_2, msg_to_bit_it_19_vnu_121_in_0, msg_to_bit_it_19_vnu_121_in_1, msg_to_bit_it_19_vnu_121_in_2, msg_to_bit_it_19_vnu_122_in_0, msg_to_bit_it_19_vnu_122_in_1, msg_to_bit_it_19_vnu_122_in_2, msg_to_bit_it_19_vnu_123_in_0, msg_to_bit_it_19_vnu_123_in_1, msg_to_bit_it_19_vnu_123_in_2, msg_to_bit_it_19_vnu_124_in_0, msg_to_bit_it_19_vnu_124_in_1, msg_to_bit_it_19_vnu_124_in_2, msg_to_bit_it_19_vnu_125_in_0, msg_to_bit_it_19_vnu_125_in_1, msg_to_bit_it_19_vnu_125_in_2, msg_to_bit_it_19_vnu_126_in_0, msg_to_bit_it_19_vnu_126_in_1, msg_to_bit_it_19_vnu_126_in_2, msg_to_bit_it_19_vnu_127_in_0, msg_to_bit_it_19_vnu_127_in_1, msg_to_bit_it_19_vnu_127_in_2, msg_to_bit_it_19_vnu_128_in_0, msg_to_bit_it_19_vnu_128_in_1, msg_to_bit_it_19_vnu_128_in_2, msg_to_bit_it_19_vnu_129_in_0, msg_to_bit_it_19_vnu_129_in_1, msg_to_bit_it_19_vnu_129_in_2, msg_to_bit_it_19_vnu_130_in_0, msg_to_bit_it_19_vnu_130_in_1, msg_to_bit_it_19_vnu_130_in_2, msg_to_bit_it_19_vnu_131_in_0, msg_to_bit_it_19_vnu_131_in_1, msg_to_bit_it_19_vnu_131_in_2, msg_to_bit_it_19_vnu_132_in_0, msg_to_bit_it_19_vnu_132_in_1, msg_to_bit_it_19_vnu_132_in_2, msg_to_bit_it_19_vnu_133_in_0, msg_to_bit_it_19_vnu_133_in_1, msg_to_bit_it_19_vnu_133_in_2, msg_to_bit_it_19_vnu_134_in_0, msg_to_bit_it_19_vnu_134_in_1, msg_to_bit_it_19_vnu_134_in_2, msg_to_bit_it_19_vnu_135_in_0, msg_to_bit_it_19_vnu_135_in_1, msg_to_bit_it_19_vnu_135_in_2, msg_to_bit_it_19_vnu_136_in_0, msg_to_bit_it_19_vnu_136_in_1, msg_to_bit_it_19_vnu_136_in_2, msg_to_bit_it_19_vnu_137_in_0, msg_to_bit_it_19_vnu_137_in_1, msg_to_bit_it_19_vnu_137_in_2, msg_to_bit_it_19_vnu_138_in_0, msg_to_bit_it_19_vnu_138_in_1, msg_to_bit_it_19_vnu_138_in_2, msg_to_bit_it_19_vnu_139_in_0, msg_to_bit_it_19_vnu_139_in_1, msg_to_bit_it_19_vnu_139_in_2, msg_to_bit_it_19_vnu_140_in_0, msg_to_bit_it_19_vnu_140_in_1, msg_to_bit_it_19_vnu_140_in_2, msg_to_bit_it_19_vnu_141_in_0, msg_to_bit_it_19_vnu_141_in_1, msg_to_bit_it_19_vnu_141_in_2, msg_to_bit_it_19_vnu_142_in_0, msg_to_bit_it_19_vnu_142_in_1, msg_to_bit_it_19_vnu_142_in_2, msg_to_bit_it_19_vnu_143_in_0, msg_to_bit_it_19_vnu_143_in_1, msg_to_bit_it_19_vnu_143_in_2, msg_to_bit_it_19_vnu_144_in_0, msg_to_bit_it_19_vnu_144_in_1, msg_to_bit_it_19_vnu_144_in_2, msg_to_bit_it_19_vnu_145_in_0, msg_to_bit_it_19_vnu_145_in_1, msg_to_bit_it_19_vnu_145_in_2, msg_to_bit_it_19_vnu_146_in_0, msg_to_bit_it_19_vnu_146_in_1, msg_to_bit_it_19_vnu_146_in_2, msg_to_bit_it_19_vnu_147_in_0, msg_to_bit_it_19_vnu_147_in_1, msg_to_bit_it_19_vnu_147_in_2, msg_to_bit_it_19_vnu_148_in_0, msg_to_bit_it_19_vnu_148_in_1, msg_to_bit_it_19_vnu_148_in_2, msg_to_bit_it_19_vnu_149_in_0, msg_to_bit_it_19_vnu_149_in_1, msg_to_bit_it_19_vnu_149_in_2, msg_to_bit_it_19_vnu_150_in_0, msg_to_bit_it_19_vnu_150_in_1, msg_to_bit_it_19_vnu_150_in_2, msg_to_bit_it_19_vnu_151_in_0, msg_to_bit_it_19_vnu_151_in_1, msg_to_bit_it_19_vnu_151_in_2, msg_to_bit_it_19_vnu_152_in_0, msg_to_bit_it_19_vnu_152_in_1, msg_to_bit_it_19_vnu_152_in_2, msg_to_bit_it_19_vnu_153_in_0, msg_to_bit_it_19_vnu_153_in_1, msg_to_bit_it_19_vnu_153_in_2, msg_to_bit_it_19_vnu_154_in_0, msg_to_bit_it_19_vnu_154_in_1, msg_to_bit_it_19_vnu_154_in_2, msg_to_bit_it_19_vnu_155_in_0, msg_to_bit_it_19_vnu_155_in_1, msg_to_bit_it_19_vnu_155_in_2, msg_to_bit_it_19_vnu_156_in_0, msg_to_bit_it_19_vnu_156_in_1, msg_to_bit_it_19_vnu_156_in_2, msg_to_bit_it_19_vnu_157_in_0, msg_to_bit_it_19_vnu_157_in_1, msg_to_bit_it_19_vnu_157_in_2, msg_to_bit_it_19_vnu_158_in_0, msg_to_bit_it_19_vnu_158_in_1, msg_to_bit_it_19_vnu_158_in_2, msg_to_bit_it_19_vnu_159_in_0, msg_to_bit_it_19_vnu_159_in_1, msg_to_bit_it_19_vnu_159_in_2, msg_to_bit_it_19_vnu_160_in_0, msg_to_bit_it_19_vnu_160_in_1, msg_to_bit_it_19_vnu_160_in_2, msg_to_bit_it_19_vnu_161_in_0, msg_to_bit_it_19_vnu_161_in_1, msg_to_bit_it_19_vnu_161_in_2, msg_to_bit_it_19_vnu_162_in_0, msg_to_bit_it_19_vnu_162_in_1, msg_to_bit_it_19_vnu_162_in_2, msg_to_bit_it_19_vnu_163_in_0, msg_to_bit_it_19_vnu_163_in_1, msg_to_bit_it_19_vnu_163_in_2, msg_to_bit_it_19_vnu_164_in_0, msg_to_bit_it_19_vnu_164_in_1, msg_to_bit_it_19_vnu_164_in_2, msg_to_bit_it_19_vnu_165_in_0, msg_to_bit_it_19_vnu_165_in_1, msg_to_bit_it_19_vnu_165_in_2, msg_to_bit_it_19_vnu_166_in_0, msg_to_bit_it_19_vnu_166_in_1, msg_to_bit_it_19_vnu_166_in_2, msg_to_bit_it_19_vnu_167_in_0, msg_to_bit_it_19_vnu_167_in_1, msg_to_bit_it_19_vnu_167_in_2, msg_to_bit_it_19_vnu_168_in_0, msg_to_bit_it_19_vnu_168_in_1, msg_to_bit_it_19_vnu_168_in_2, msg_to_bit_it_19_vnu_169_in_0, msg_to_bit_it_19_vnu_169_in_1, msg_to_bit_it_19_vnu_169_in_2, msg_to_bit_it_19_vnu_170_in_0, msg_to_bit_it_19_vnu_170_in_1, msg_to_bit_it_19_vnu_170_in_2, msg_to_bit_it_19_vnu_171_in_0, msg_to_bit_it_19_vnu_171_in_1, msg_to_bit_it_19_vnu_171_in_2, msg_to_bit_it_19_vnu_172_in_0, msg_to_bit_it_19_vnu_172_in_1, msg_to_bit_it_19_vnu_172_in_2, msg_to_bit_it_19_vnu_173_in_0, msg_to_bit_it_19_vnu_173_in_1, msg_to_bit_it_19_vnu_173_in_2, msg_to_bit_it_19_vnu_174_in_0, msg_to_bit_it_19_vnu_174_in_1, msg_to_bit_it_19_vnu_174_in_2, msg_to_bit_it_19_vnu_175_in_0, msg_to_bit_it_19_vnu_175_in_1, msg_to_bit_it_19_vnu_175_in_2, msg_to_bit_it_19_vnu_176_in_0, msg_to_bit_it_19_vnu_176_in_1, msg_to_bit_it_19_vnu_176_in_2, msg_to_bit_it_19_vnu_177_in_0, msg_to_bit_it_19_vnu_177_in_1, msg_to_bit_it_19_vnu_177_in_2, msg_to_bit_it_19_vnu_178_in_0, msg_to_bit_it_19_vnu_178_in_1, msg_to_bit_it_19_vnu_178_in_2, msg_to_bit_it_19_vnu_179_in_0, msg_to_bit_it_19_vnu_179_in_1, msg_to_bit_it_19_vnu_179_in_2, msg_to_bit_it_19_vnu_180_in_0, msg_to_bit_it_19_vnu_180_in_1, msg_to_bit_it_19_vnu_180_in_2, msg_to_bit_it_19_vnu_181_in_0, msg_to_bit_it_19_vnu_181_in_1, msg_to_bit_it_19_vnu_181_in_2, msg_to_bit_it_19_vnu_182_in_0, msg_to_bit_it_19_vnu_182_in_1, msg_to_bit_it_19_vnu_182_in_2, msg_to_bit_it_19_vnu_183_in_0, msg_to_bit_it_19_vnu_183_in_1, msg_to_bit_it_19_vnu_183_in_2, msg_to_bit_it_19_vnu_184_in_0, msg_to_bit_it_19_vnu_184_in_1, msg_to_bit_it_19_vnu_184_in_2, msg_to_bit_it_19_vnu_185_in_0, msg_to_bit_it_19_vnu_185_in_1, msg_to_bit_it_19_vnu_185_in_2, msg_to_bit_it_19_vnu_186_in_0, msg_to_bit_it_19_vnu_186_in_1, msg_to_bit_it_19_vnu_186_in_2, msg_to_bit_it_19_vnu_187_in_0, msg_to_bit_it_19_vnu_187_in_1, msg_to_bit_it_19_vnu_187_in_2, msg_to_bit_it_19_vnu_188_in_0, msg_to_bit_it_19_vnu_188_in_1, msg_to_bit_it_19_vnu_188_in_2, msg_to_bit_it_19_vnu_189_in_0, msg_to_bit_it_19_vnu_189_in_1, msg_to_bit_it_19_vnu_189_in_2, msg_to_bit_it_19_vnu_190_in_0, msg_to_bit_it_19_vnu_190_in_1, msg_to_bit_it_19_vnu_190_in_2, msg_to_bit_it_19_vnu_191_in_0, msg_to_bit_it_19_vnu_191_in_1, msg_to_bit_it_19_vnu_191_in_2, msg_to_bit_it_19_vnu_192_in_0, msg_to_bit_it_19_vnu_192_in_1, msg_to_bit_it_19_vnu_192_in_2, msg_to_bit_it_19_vnu_193_in_0, msg_to_bit_it_19_vnu_193_in_1, msg_to_bit_it_19_vnu_193_in_2, msg_to_bit_it_19_vnu_194_in_0, msg_to_bit_it_19_vnu_194_in_1, msg_to_bit_it_19_vnu_194_in_2, msg_to_bit_it_19_vnu_195_in_0, msg_to_bit_it_19_vnu_195_in_1, msg_to_bit_it_19_vnu_195_in_2, msg_to_bit_it_19_vnu_196_in_0, msg_to_bit_it_19_vnu_196_in_1, msg_to_bit_it_19_vnu_196_in_2, msg_to_bit_it_19_vnu_197_in_0, msg_to_bit_it_19_vnu_197_in_1, msg_to_bit_it_19_vnu_197_in_2;
//reg decode_in_en;
//wire clk;
//always @(data_in_en) begin
//	decode_in_en = 1;
//end

wire cnu_over, vnu_over;
reg decode_en, vnu_en, cnu_en, get_output;

always @(posedge clk) begin
	if(~rst) begin
		decode_en = 0;
		vnu_en = 0;
		cnu_en = 0;
	end
	else begin
		decode_en = 1;	
		vnu_en = 1;
		//cnu_en = 1;
	end
end

always @(vnu_over) begin
	if(vnu_over == 1)
		cnu_en = 1;
end
//for other iterations continue
always @(cnu_over) begin
	if(cnu_over == 1) begin
		get_output = 1;
	end
end




vnu_1 variable_node_0_0(data_0, msg_to_check_it_0_cnu_31_in_0, msg_to_check_it_0_cnu_62_in_0, msg_to_check_it_0_cnu_93_in_0);
vnu_1 variable_node_1_0(data_1, msg_to_check_it_0_cnu_32_in_0, msg_to_check_it_0_cnu_63_in_0, msg_to_check_it_0_cnu_94_in_0);
vnu_1 variable_node_2_0(data_2, msg_to_check_it_0_cnu_0_in_0, msg_to_check_it_0_cnu_64_in_0, msg_to_check_it_0_cnu_95_in_0);
vnu_1 variable_node_3_0(data_3, msg_to_check_it_0_cnu_1_in_0, msg_to_check_it_0_cnu_65_in_0, msg_to_check_it_0_cnu_96_in_0);
vnu_1 variable_node_4_0(data_4, msg_to_check_it_0_cnu_2_in_0, msg_to_check_it_0_cnu_33_in_0, msg_to_check_it_0_cnu_97_in_0);
vnu_1 variable_node_5_0(data_5, msg_to_check_it_0_cnu_3_in_0, msg_to_check_it_0_cnu_34_in_0, msg_to_check_it_0_cnu_98_in_0);
vnu_1 variable_node_6_0(data_6, msg_to_check_it_0_cnu_4_in_0, msg_to_check_it_0_cnu_35_in_0, msg_to_check_it_0_cnu_66_in_0);
vnu_1 variable_node_7_0(data_7, msg_to_check_it_0_cnu_5_in_0, msg_to_check_it_0_cnu_36_in_0, msg_to_check_it_0_cnu_67_in_0);
vnu_1 variable_node_8_0(data_8, msg_to_check_it_0_cnu_6_in_0, msg_to_check_it_0_cnu_37_in_0, msg_to_check_it_0_cnu_68_in_0);
vnu_1 variable_node_9_0(data_9, msg_to_check_it_0_cnu_7_in_0, msg_to_check_it_0_cnu_38_in_0, msg_to_check_it_0_cnu_69_in_0);
vnu_1 variable_node_10_0(data_10, msg_to_check_it_0_cnu_8_in_0, msg_to_check_it_0_cnu_39_in_0, msg_to_check_it_0_cnu_70_in_0);
vnu_1 variable_node_11_0(data_11, msg_to_check_it_0_cnu_9_in_0, msg_to_check_it_0_cnu_40_in_0, msg_to_check_it_0_cnu_71_in_0);
vnu_1 variable_node_12_0(data_12, msg_to_check_it_0_cnu_10_in_0, msg_to_check_it_0_cnu_41_in_0, msg_to_check_it_0_cnu_72_in_0);
vnu_1 variable_node_13_0(data_13, msg_to_check_it_0_cnu_11_in_0, msg_to_check_it_0_cnu_42_in_0, msg_to_check_it_0_cnu_73_in_0);
vnu_1 variable_node_14_0(data_14, msg_to_check_it_0_cnu_12_in_0, msg_to_check_it_0_cnu_43_in_0, msg_to_check_it_0_cnu_74_in_0);
vnu_1 variable_node_15_0(data_15, msg_to_check_it_0_cnu_13_in_0, msg_to_check_it_0_cnu_44_in_0, msg_to_check_it_0_cnu_75_in_0);
vnu_1 variable_node_16_0(data_16, msg_to_check_it_0_cnu_14_in_0, msg_to_check_it_0_cnu_45_in_0, msg_to_check_it_0_cnu_76_in_0);
vnu_1 variable_node_17_0(data_17, msg_to_check_it_0_cnu_15_in_0, msg_to_check_it_0_cnu_46_in_0, msg_to_check_it_0_cnu_77_in_0);
vnu_1 variable_node_18_0(data_18, msg_to_check_it_0_cnu_16_in_0, msg_to_check_it_0_cnu_47_in_0, msg_to_check_it_0_cnu_78_in_0);
vnu_1 variable_node_19_0(data_19, msg_to_check_it_0_cnu_17_in_0, msg_to_check_it_0_cnu_48_in_0, msg_to_check_it_0_cnu_79_in_0);
vnu_1 variable_node_20_0(data_20, msg_to_check_it_0_cnu_18_in_0, msg_to_check_it_0_cnu_49_in_0, msg_to_check_it_0_cnu_80_in_0);
vnu_1 variable_node_21_0(data_21, msg_to_check_it_0_cnu_19_in_0, msg_to_check_it_0_cnu_50_in_0, msg_to_check_it_0_cnu_81_in_0);
vnu_1 variable_node_22_0(data_22, msg_to_check_it_0_cnu_20_in_0, msg_to_check_it_0_cnu_51_in_0, msg_to_check_it_0_cnu_82_in_0);
vnu_1 variable_node_23_0(data_23, msg_to_check_it_0_cnu_21_in_0, msg_to_check_it_0_cnu_52_in_0, msg_to_check_it_0_cnu_83_in_0);
vnu_1 variable_node_24_0(data_24, msg_to_check_it_0_cnu_22_in_0, msg_to_check_it_0_cnu_53_in_0, msg_to_check_it_0_cnu_84_in_0);
vnu_1 variable_node_25_0(data_25, msg_to_check_it_0_cnu_23_in_0, msg_to_check_it_0_cnu_54_in_0, msg_to_check_it_0_cnu_85_in_0);
vnu_1 variable_node_26_0(data_26, msg_to_check_it_0_cnu_24_in_0, msg_to_check_it_0_cnu_55_in_0, msg_to_check_it_0_cnu_86_in_0);
vnu_1 variable_node_27_0(data_27, msg_to_check_it_0_cnu_25_in_0, msg_to_check_it_0_cnu_56_in_0, msg_to_check_it_0_cnu_87_in_0);
vnu_1 variable_node_28_0(data_28, msg_to_check_it_0_cnu_26_in_0, msg_to_check_it_0_cnu_57_in_0, msg_to_check_it_0_cnu_88_in_0);
vnu_1 variable_node_29_0(data_29, msg_to_check_it_0_cnu_27_in_0, msg_to_check_it_0_cnu_58_in_0, msg_to_check_it_0_cnu_89_in_0);
vnu_1 variable_node_30_0(data_30, msg_to_check_it_0_cnu_28_in_0, msg_to_check_it_0_cnu_59_in_0, msg_to_check_it_0_cnu_90_in_0);
vnu_1 variable_node_31_0(data_31, msg_to_check_it_0_cnu_29_in_0, msg_to_check_it_0_cnu_60_in_0, msg_to_check_it_0_cnu_91_in_0);
vnu_1 variable_node_32_0(data_32, msg_to_check_it_0_cnu_30_in_0, msg_to_check_it_0_cnu_61_in_0, msg_to_check_it_0_cnu_92_in_0);
vnu_1 variable_node_33_0(data_33, msg_to_check_it_0_cnu_30_in_1, msg_to_check_it_0_cnu_61_in_1, msg_to_check_it_0_cnu_91_in_1);
vnu_1 variable_node_34_0(data_34, msg_to_check_it_0_cnu_31_in_1, msg_to_check_it_0_cnu_62_in_1, msg_to_check_it_0_cnu_92_in_1);
vnu_1 variable_node_35_0(data_35, msg_to_check_it_0_cnu_32_in_1, msg_to_check_it_0_cnu_63_in_1, msg_to_check_it_0_cnu_93_in_1);
vnu_1 variable_node_36_0(data_36, msg_to_check_it_0_cnu_0_in_1, msg_to_check_it_0_cnu_64_in_1, msg_to_check_it_0_cnu_94_in_1);
vnu_1 variable_node_37_0(data_37, msg_to_check_it_0_cnu_1_in_1, msg_to_check_it_0_cnu_65_in_1, msg_to_check_it_0_cnu_95_in_1);
vnu_1 variable_node_38_0(data_38, msg_to_check_it_0_cnu_2_in_1, msg_to_check_it_0_cnu_33_in_1, msg_to_check_it_0_cnu_96_in_1);
vnu_1 variable_node_39_0(data_39, msg_to_check_it_0_cnu_3_in_1, msg_to_check_it_0_cnu_34_in_1, msg_to_check_it_0_cnu_97_in_1);
vnu_1 variable_node_40_0(data_40, msg_to_check_it_0_cnu_4_in_1, msg_to_check_it_0_cnu_35_in_1, msg_to_check_it_0_cnu_98_in_1);
vnu_1 variable_node_41_0(data_41, msg_to_check_it_0_cnu_5_in_1, msg_to_check_it_0_cnu_36_in_1, msg_to_check_it_0_cnu_66_in_1);
vnu_1 variable_node_42_0(data_42, msg_to_check_it_0_cnu_6_in_1, msg_to_check_it_0_cnu_37_in_1, msg_to_check_it_0_cnu_67_in_1);
vnu_1 variable_node_43_0(data_43, msg_to_check_it_0_cnu_7_in_1, msg_to_check_it_0_cnu_38_in_1, msg_to_check_it_0_cnu_68_in_1);
vnu_1 variable_node_44_0(data_44, msg_to_check_it_0_cnu_8_in_1, msg_to_check_it_0_cnu_39_in_1, msg_to_check_it_0_cnu_69_in_1);
vnu_1 variable_node_45_0(data_45, msg_to_check_it_0_cnu_9_in_1, msg_to_check_it_0_cnu_40_in_1, msg_to_check_it_0_cnu_70_in_1);
vnu_1 variable_node_46_0(data_46, msg_to_check_it_0_cnu_10_in_1, msg_to_check_it_0_cnu_41_in_1, msg_to_check_it_0_cnu_71_in_1);
vnu_1 variable_node_47_0(data_47, msg_to_check_it_0_cnu_11_in_1, msg_to_check_it_0_cnu_42_in_1, msg_to_check_it_0_cnu_72_in_1);
vnu_1 variable_node_48_0(data_48, msg_to_check_it_0_cnu_12_in_1, msg_to_check_it_0_cnu_43_in_1, msg_to_check_it_0_cnu_73_in_1);
vnu_1 variable_node_49_0(data_49, msg_to_check_it_0_cnu_13_in_1, msg_to_check_it_0_cnu_44_in_1, msg_to_check_it_0_cnu_74_in_1);
vnu_1 variable_node_50_0(data_50, msg_to_check_it_0_cnu_14_in_1, msg_to_check_it_0_cnu_45_in_1, msg_to_check_it_0_cnu_75_in_1);
vnu_1 variable_node_51_0(data_51, msg_to_check_it_0_cnu_15_in_1, msg_to_check_it_0_cnu_46_in_1, msg_to_check_it_0_cnu_76_in_1);
vnu_1 variable_node_52_0(data_52, msg_to_check_it_0_cnu_16_in_1, msg_to_check_it_0_cnu_47_in_1, msg_to_check_it_0_cnu_77_in_1);
vnu_1 variable_node_53_0(data_53, msg_to_check_it_0_cnu_17_in_1, msg_to_check_it_0_cnu_48_in_1, msg_to_check_it_0_cnu_78_in_1);
vnu_1 variable_node_54_0(data_54, msg_to_check_it_0_cnu_18_in_1, msg_to_check_it_0_cnu_49_in_1, msg_to_check_it_0_cnu_79_in_1);
vnu_1 variable_node_55_0(data_55, msg_to_check_it_0_cnu_19_in_1, msg_to_check_it_0_cnu_50_in_1, msg_to_check_it_0_cnu_80_in_1);
vnu_1 variable_node_56_0(data_56, msg_to_check_it_0_cnu_20_in_1, msg_to_check_it_0_cnu_51_in_1, msg_to_check_it_0_cnu_81_in_1);
vnu_1 variable_node_57_0(data_57, msg_to_check_it_0_cnu_21_in_1, msg_to_check_it_0_cnu_52_in_1, msg_to_check_it_0_cnu_82_in_1);
vnu_1 variable_node_58_0(data_58, msg_to_check_it_0_cnu_22_in_1, msg_to_check_it_0_cnu_53_in_1, msg_to_check_it_0_cnu_83_in_1);
vnu_1 variable_node_59_0(data_59, msg_to_check_it_0_cnu_23_in_1, msg_to_check_it_0_cnu_54_in_1, msg_to_check_it_0_cnu_84_in_1);
vnu_1 variable_node_60_0(data_60, msg_to_check_it_0_cnu_24_in_1, msg_to_check_it_0_cnu_55_in_1, msg_to_check_it_0_cnu_85_in_1);
vnu_1 variable_node_61_0(data_61, msg_to_check_it_0_cnu_25_in_1, msg_to_check_it_0_cnu_56_in_1, msg_to_check_it_0_cnu_86_in_1);
vnu_1 variable_node_62_0(data_62, msg_to_check_it_0_cnu_26_in_1, msg_to_check_it_0_cnu_57_in_1, msg_to_check_it_0_cnu_87_in_1);
vnu_1 variable_node_63_0(data_63, msg_to_check_it_0_cnu_27_in_1, msg_to_check_it_0_cnu_58_in_1, msg_to_check_it_0_cnu_88_in_1);
vnu_1 variable_node_64_0(data_64, msg_to_check_it_0_cnu_28_in_1, msg_to_check_it_0_cnu_59_in_1, msg_to_check_it_0_cnu_89_in_1);
vnu_1 variable_node_65_0(data_65, msg_to_check_it_0_cnu_29_in_1, msg_to_check_it_0_cnu_60_in_1, msg_to_check_it_0_cnu_90_in_1);
vnu_1 variable_node_66_0(data_66, msg_to_check_it_0_cnu_26_in_2, msg_to_check_it_0_cnu_55_in_2, msg_to_check_it_0_cnu_85_in_2);
vnu_1 variable_node_67_0(data_67, msg_to_check_it_0_cnu_27_in_2, msg_to_check_it_0_cnu_56_in_2, msg_to_check_it_0_cnu_86_in_2);
vnu_1 variable_node_68_0(data_68, msg_to_check_it_0_cnu_28_in_2, msg_to_check_it_0_cnu_57_in_2, msg_to_check_it_0_cnu_87_in_2);
vnu_1 variable_node_69_0(data_69, msg_to_check_it_0_cnu_29_in_2, msg_to_check_it_0_cnu_58_in_2, msg_to_check_it_0_cnu_88_in_2);
vnu_1 variable_node_70_0(data_70, msg_to_check_it_0_cnu_30_in_2, msg_to_check_it_0_cnu_59_in_2, msg_to_check_it_0_cnu_89_in_2);
vnu_1 variable_node_71_0(data_71, msg_to_check_it_0_cnu_31_in_2, msg_to_check_it_0_cnu_60_in_2, msg_to_check_it_0_cnu_90_in_2);
vnu_1 variable_node_72_0(data_72, msg_to_check_it_0_cnu_32_in_2, msg_to_check_it_0_cnu_61_in_2, msg_to_check_it_0_cnu_91_in_2);
vnu_1 variable_node_73_0(data_73, msg_to_check_it_0_cnu_0_in_2, msg_to_check_it_0_cnu_62_in_2, msg_to_check_it_0_cnu_92_in_2);
vnu_1 variable_node_74_0(data_74, msg_to_check_it_0_cnu_1_in_2, msg_to_check_it_0_cnu_63_in_2, msg_to_check_it_0_cnu_93_in_2);
vnu_1 variable_node_75_0(data_75, msg_to_check_it_0_cnu_2_in_2, msg_to_check_it_0_cnu_64_in_2, msg_to_check_it_0_cnu_94_in_2);
vnu_1 variable_node_76_0(data_76, msg_to_check_it_0_cnu_3_in_2, msg_to_check_it_0_cnu_65_in_2, msg_to_check_it_0_cnu_95_in_2);
vnu_1 variable_node_77_0(data_77, msg_to_check_it_0_cnu_4_in_2, msg_to_check_it_0_cnu_33_in_2, msg_to_check_it_0_cnu_96_in_2);
vnu_1 variable_node_78_0(data_78, msg_to_check_it_0_cnu_5_in_2, msg_to_check_it_0_cnu_34_in_2, msg_to_check_it_0_cnu_97_in_2);
vnu_1 variable_node_79_0(data_79, msg_to_check_it_0_cnu_6_in_2, msg_to_check_it_0_cnu_35_in_2, msg_to_check_it_0_cnu_98_in_2);
vnu_1 variable_node_80_0(data_80, msg_to_check_it_0_cnu_7_in_2, msg_to_check_it_0_cnu_36_in_2, msg_to_check_it_0_cnu_66_in_2);
vnu_1 variable_node_81_0(data_81, msg_to_check_it_0_cnu_8_in_2, msg_to_check_it_0_cnu_37_in_2, msg_to_check_it_0_cnu_67_in_2);
vnu_1 variable_node_82_0(data_82, msg_to_check_it_0_cnu_9_in_2, msg_to_check_it_0_cnu_38_in_2, msg_to_check_it_0_cnu_68_in_2);
vnu_1 variable_node_83_0(data_83, msg_to_check_it_0_cnu_10_in_2, msg_to_check_it_0_cnu_39_in_2, msg_to_check_it_0_cnu_69_in_2);
vnu_1 variable_node_84_0(data_84, msg_to_check_it_0_cnu_11_in_2, msg_to_check_it_0_cnu_40_in_2, msg_to_check_it_0_cnu_70_in_2);
vnu_1 variable_node_85_0(data_85, msg_to_check_it_0_cnu_12_in_2, msg_to_check_it_0_cnu_41_in_2, msg_to_check_it_0_cnu_71_in_2);
vnu_1 variable_node_86_0(data_86, msg_to_check_it_0_cnu_13_in_2, msg_to_check_it_0_cnu_42_in_2, msg_to_check_it_0_cnu_72_in_2);
vnu_1 variable_node_87_0(data_87, msg_to_check_it_0_cnu_14_in_2, msg_to_check_it_0_cnu_43_in_2, msg_to_check_it_0_cnu_73_in_2);
vnu_1 variable_node_88_0(data_88, msg_to_check_it_0_cnu_15_in_2, msg_to_check_it_0_cnu_44_in_2, msg_to_check_it_0_cnu_74_in_2);
vnu_1 variable_node_89_0(data_89, msg_to_check_it_0_cnu_16_in_2, msg_to_check_it_0_cnu_45_in_2, msg_to_check_it_0_cnu_75_in_2);
vnu_1 variable_node_90_0(data_90, msg_to_check_it_0_cnu_17_in_2, msg_to_check_it_0_cnu_46_in_2, msg_to_check_it_0_cnu_76_in_2);
vnu_1 variable_node_91_0(data_91, msg_to_check_it_0_cnu_18_in_2, msg_to_check_it_0_cnu_47_in_2, msg_to_check_it_0_cnu_77_in_2);
vnu_1 variable_node_92_0(data_92, msg_to_check_it_0_cnu_19_in_2, msg_to_check_it_0_cnu_48_in_2, msg_to_check_it_0_cnu_78_in_2);
vnu_1 variable_node_93_0(data_93, msg_to_check_it_0_cnu_20_in_2, msg_to_check_it_0_cnu_49_in_2, msg_to_check_it_0_cnu_79_in_2);
vnu_1 variable_node_94_0(data_94, msg_to_check_it_0_cnu_21_in_2, msg_to_check_it_0_cnu_50_in_2, msg_to_check_it_0_cnu_80_in_2);
vnu_1 variable_node_95_0(data_95, msg_to_check_it_0_cnu_22_in_2, msg_to_check_it_0_cnu_51_in_2, msg_to_check_it_0_cnu_81_in_2);
vnu_1 variable_node_96_0(data_96, msg_to_check_it_0_cnu_23_in_2, msg_to_check_it_0_cnu_52_in_2, msg_to_check_it_0_cnu_82_in_2);
vnu_1 variable_node_97_0(data_97, msg_to_check_it_0_cnu_24_in_2, msg_to_check_it_0_cnu_53_in_2, msg_to_check_it_0_cnu_83_in_2);
vnu_1 variable_node_98_0(data_98, msg_to_check_it_0_cnu_25_in_2, msg_to_check_it_0_cnu_54_in_2, msg_to_check_it_0_cnu_84_in_2);
vnu_1 variable_node_99_0(data_99, msg_to_check_it_0_cnu_24_in_3, msg_to_check_it_0_cnu_54_in_3, msg_to_check_it_0_cnu_80_in_3);
vnu_1 variable_node_100_0(data_100, msg_to_check_it_0_cnu_25_in_3, msg_to_check_it_0_cnu_55_in_3, msg_to_check_it_0_cnu_81_in_3);
vnu_1 variable_node_101_0(data_101, msg_to_check_it_0_cnu_26_in_3, msg_to_check_it_0_cnu_56_in_3, msg_to_check_it_0_cnu_82_in_3);
vnu_1 variable_node_102_0(data_102, msg_to_check_it_0_cnu_27_in_3, msg_to_check_it_0_cnu_57_in_3, msg_to_check_it_0_cnu_83_in_3);
vnu_1 variable_node_103_0(data_103, msg_to_check_it_0_cnu_28_in_3, msg_to_check_it_0_cnu_58_in_3, msg_to_check_it_0_cnu_84_in_3);
vnu_1 variable_node_104_0(data_104, msg_to_check_it_0_cnu_29_in_3, msg_to_check_it_0_cnu_59_in_3, msg_to_check_it_0_cnu_85_in_3);
vnu_1 variable_node_105_0(data_105, msg_to_check_it_0_cnu_30_in_3, msg_to_check_it_0_cnu_60_in_3, msg_to_check_it_0_cnu_86_in_3);
vnu_1 variable_node_106_0(data_106, msg_to_check_it_0_cnu_31_in_3, msg_to_check_it_0_cnu_61_in_3, msg_to_check_it_0_cnu_87_in_3);
vnu_1 variable_node_107_0(data_107, msg_to_check_it_0_cnu_32_in_3, msg_to_check_it_0_cnu_62_in_3, msg_to_check_it_0_cnu_88_in_3);
vnu_1 variable_node_108_0(data_108, msg_to_check_it_0_cnu_0_in_3, msg_to_check_it_0_cnu_63_in_3, msg_to_check_it_0_cnu_89_in_3);
vnu_1 variable_node_109_0(data_109, msg_to_check_it_0_cnu_1_in_3, msg_to_check_it_0_cnu_64_in_3, msg_to_check_it_0_cnu_90_in_3);
vnu_1 variable_node_110_0(data_110, msg_to_check_it_0_cnu_2_in_3, msg_to_check_it_0_cnu_65_in_3, msg_to_check_it_0_cnu_91_in_3);
vnu_1 variable_node_111_0(data_111, msg_to_check_it_0_cnu_3_in_3, msg_to_check_it_0_cnu_33_in_3, msg_to_check_it_0_cnu_92_in_3);
vnu_1 variable_node_112_0(data_112, msg_to_check_it_0_cnu_4_in_3, msg_to_check_it_0_cnu_34_in_3, msg_to_check_it_0_cnu_93_in_3);
vnu_1 variable_node_113_0(data_113, msg_to_check_it_0_cnu_5_in_3, msg_to_check_it_0_cnu_35_in_3, msg_to_check_it_0_cnu_94_in_3);
vnu_1 variable_node_114_0(data_114, msg_to_check_it_0_cnu_6_in_3, msg_to_check_it_0_cnu_36_in_3, msg_to_check_it_0_cnu_95_in_3);
vnu_1 variable_node_115_0(data_115, msg_to_check_it_0_cnu_7_in_3, msg_to_check_it_0_cnu_37_in_3, msg_to_check_it_0_cnu_96_in_3);
vnu_1 variable_node_116_0(data_116, msg_to_check_it_0_cnu_8_in_3, msg_to_check_it_0_cnu_38_in_3, msg_to_check_it_0_cnu_97_in_3);
vnu_1 variable_node_117_0(data_117, msg_to_check_it_0_cnu_9_in_3, msg_to_check_it_0_cnu_39_in_3, msg_to_check_it_0_cnu_98_in_3);
vnu_1 variable_node_118_0(data_118, msg_to_check_it_0_cnu_10_in_3, msg_to_check_it_0_cnu_40_in_3, msg_to_check_it_0_cnu_66_in_3);
vnu_1 variable_node_119_0(data_119, msg_to_check_it_0_cnu_11_in_3, msg_to_check_it_0_cnu_41_in_3, msg_to_check_it_0_cnu_67_in_3);
vnu_1 variable_node_120_0(data_120, msg_to_check_it_0_cnu_12_in_3, msg_to_check_it_0_cnu_42_in_3, msg_to_check_it_0_cnu_68_in_3);
vnu_1 variable_node_121_0(data_121, msg_to_check_it_0_cnu_13_in_3, msg_to_check_it_0_cnu_43_in_3, msg_to_check_it_0_cnu_69_in_3);
vnu_1 variable_node_122_0(data_122, msg_to_check_it_0_cnu_14_in_3, msg_to_check_it_0_cnu_44_in_3, msg_to_check_it_0_cnu_70_in_3);
vnu_1 variable_node_123_0(data_123, msg_to_check_it_0_cnu_15_in_3, msg_to_check_it_0_cnu_45_in_3, msg_to_check_it_0_cnu_71_in_3);
vnu_1 variable_node_124_0(data_124, msg_to_check_it_0_cnu_16_in_3, msg_to_check_it_0_cnu_46_in_3, msg_to_check_it_0_cnu_72_in_3);
vnu_1 variable_node_125_0(data_125, msg_to_check_it_0_cnu_17_in_3, msg_to_check_it_0_cnu_47_in_3, msg_to_check_it_0_cnu_73_in_3);
vnu_1 variable_node_126_0(data_126, msg_to_check_it_0_cnu_18_in_3, msg_to_check_it_0_cnu_48_in_3, msg_to_check_it_0_cnu_74_in_3);
vnu_1 variable_node_127_0(data_127, msg_to_check_it_0_cnu_19_in_3, msg_to_check_it_0_cnu_49_in_3, msg_to_check_it_0_cnu_75_in_3);
vnu_1 variable_node_128_0(data_128, msg_to_check_it_0_cnu_20_in_3, msg_to_check_it_0_cnu_50_in_3, msg_to_check_it_0_cnu_76_in_3);
vnu_1 variable_node_129_0(data_129, msg_to_check_it_0_cnu_21_in_3, msg_to_check_it_0_cnu_51_in_3, msg_to_check_it_0_cnu_77_in_3);
vnu_1 variable_node_130_0(data_130, msg_to_check_it_0_cnu_22_in_3, msg_to_check_it_0_cnu_52_in_3, msg_to_check_it_0_cnu_78_in_3);
vnu_1 variable_node_131_0(data_131, msg_to_check_it_0_cnu_23_in_3, msg_to_check_it_0_cnu_53_in_3, msg_to_check_it_0_cnu_79_in_3);
vnu_1 variable_node_132_0(data_132, msg_to_check_it_0_cnu_18_in_4, msg_to_check_it_0_cnu_43_in_4, msg_to_check_it_0_cnu_72_in_4);
vnu_1 variable_node_133_0(data_133, msg_to_check_it_0_cnu_19_in_4, msg_to_check_it_0_cnu_44_in_4, msg_to_check_it_0_cnu_73_in_4);
vnu_1 variable_node_134_0(data_134, msg_to_check_it_0_cnu_20_in_4, msg_to_check_it_0_cnu_45_in_4, msg_to_check_it_0_cnu_74_in_4);
vnu_1 variable_node_135_0(data_135, msg_to_check_it_0_cnu_21_in_4, msg_to_check_it_0_cnu_46_in_4, msg_to_check_it_0_cnu_75_in_4);
vnu_1 variable_node_136_0(data_136, msg_to_check_it_0_cnu_22_in_4, msg_to_check_it_0_cnu_47_in_4, msg_to_check_it_0_cnu_76_in_4);
vnu_1 variable_node_137_0(data_137, msg_to_check_it_0_cnu_23_in_4, msg_to_check_it_0_cnu_48_in_4, msg_to_check_it_0_cnu_77_in_4);
vnu_1 variable_node_138_0(data_138, msg_to_check_it_0_cnu_24_in_4, msg_to_check_it_0_cnu_49_in_4, msg_to_check_it_0_cnu_78_in_4);
vnu_1 variable_node_139_0(data_139, msg_to_check_it_0_cnu_25_in_4, msg_to_check_it_0_cnu_50_in_4, msg_to_check_it_0_cnu_79_in_4);
vnu_1 variable_node_140_0(data_140, msg_to_check_it_0_cnu_26_in_4, msg_to_check_it_0_cnu_51_in_4, msg_to_check_it_0_cnu_80_in_4);
vnu_1 variable_node_141_0(data_141, msg_to_check_it_0_cnu_27_in_4, msg_to_check_it_0_cnu_52_in_4, msg_to_check_it_0_cnu_81_in_4);
vnu_1 variable_node_142_0(data_142, msg_to_check_it_0_cnu_28_in_4, msg_to_check_it_0_cnu_53_in_4, msg_to_check_it_0_cnu_82_in_4);
vnu_1 variable_node_143_0(data_143, msg_to_check_it_0_cnu_29_in_4, msg_to_check_it_0_cnu_54_in_4, msg_to_check_it_0_cnu_83_in_4);
vnu_1 variable_node_144_0(data_144, msg_to_check_it_0_cnu_30_in_4, msg_to_check_it_0_cnu_55_in_4, msg_to_check_it_0_cnu_84_in_4);
vnu_1 variable_node_145_0(data_145, msg_to_check_it_0_cnu_31_in_4, msg_to_check_it_0_cnu_56_in_4, msg_to_check_it_0_cnu_85_in_4);
vnu_1 variable_node_146_0(data_146, msg_to_check_it_0_cnu_32_in_4, msg_to_check_it_0_cnu_57_in_4, msg_to_check_it_0_cnu_86_in_4);
vnu_1 variable_node_147_0(data_147, msg_to_check_it_0_cnu_0_in_4, msg_to_check_it_0_cnu_58_in_4, msg_to_check_it_0_cnu_87_in_4);
vnu_1 variable_node_148_0(data_148, msg_to_check_it_0_cnu_1_in_4, msg_to_check_it_0_cnu_59_in_4, msg_to_check_it_0_cnu_88_in_4);
vnu_1 variable_node_149_0(data_149, msg_to_check_it_0_cnu_2_in_4, msg_to_check_it_0_cnu_60_in_4, msg_to_check_it_0_cnu_89_in_4);
vnu_1 variable_node_150_0(data_150, msg_to_check_it_0_cnu_3_in_4, msg_to_check_it_0_cnu_61_in_4, msg_to_check_it_0_cnu_90_in_4);
vnu_1 variable_node_151_0(data_151, msg_to_check_it_0_cnu_4_in_4, msg_to_check_it_0_cnu_62_in_4, msg_to_check_it_0_cnu_91_in_4);
vnu_1 variable_node_152_0(data_152, msg_to_check_it_0_cnu_5_in_4, msg_to_check_it_0_cnu_63_in_4, msg_to_check_it_0_cnu_92_in_4);
vnu_1 variable_node_153_0(data_153, msg_to_check_it_0_cnu_6_in_4, msg_to_check_it_0_cnu_64_in_4, msg_to_check_it_0_cnu_93_in_4);
vnu_1 variable_node_154_0(data_154, msg_to_check_it_0_cnu_7_in_4, msg_to_check_it_0_cnu_65_in_4, msg_to_check_it_0_cnu_94_in_4);
vnu_1 variable_node_155_0(data_155, msg_to_check_it_0_cnu_8_in_4, msg_to_check_it_0_cnu_33_in_4, msg_to_check_it_0_cnu_95_in_4);
vnu_1 variable_node_156_0(data_156, msg_to_check_it_0_cnu_9_in_4, msg_to_check_it_0_cnu_34_in_4, msg_to_check_it_0_cnu_96_in_4);
vnu_1 variable_node_157_0(data_157, msg_to_check_it_0_cnu_10_in_4, msg_to_check_it_0_cnu_35_in_4, msg_to_check_it_0_cnu_97_in_4);
vnu_1 variable_node_158_0(data_158, msg_to_check_it_0_cnu_11_in_4, msg_to_check_it_0_cnu_36_in_4, msg_to_check_it_0_cnu_98_in_4);
vnu_1 variable_node_159_0(data_159, msg_to_check_it_0_cnu_12_in_4, msg_to_check_it_0_cnu_37_in_4, msg_to_check_it_0_cnu_66_in_4);
vnu_1 variable_node_160_0(data_160, msg_to_check_it_0_cnu_13_in_4, msg_to_check_it_0_cnu_38_in_4, msg_to_check_it_0_cnu_67_in_4);
vnu_1 variable_node_161_0(data_161, msg_to_check_it_0_cnu_14_in_4, msg_to_check_it_0_cnu_39_in_4, msg_to_check_it_0_cnu_68_in_4);
vnu_1 variable_node_162_0(data_162, msg_to_check_it_0_cnu_15_in_4, msg_to_check_it_0_cnu_40_in_4, msg_to_check_it_0_cnu_69_in_4);
vnu_1 variable_node_163_0(data_163, msg_to_check_it_0_cnu_16_in_4, msg_to_check_it_0_cnu_41_in_4, msg_to_check_it_0_cnu_70_in_4);
vnu_1 variable_node_164_0(data_164, msg_to_check_it_0_cnu_17_in_4, msg_to_check_it_0_cnu_42_in_4, msg_to_check_it_0_cnu_71_in_4);
vnu_1 variable_node_165_0(data_165, msg_to_check_it_0_cnu_13_in_5, msg_to_check_it_0_cnu_41_in_5, msg_to_check_it_0_cnu_69_in_5);
vnu_1 variable_node_166_0(data_166, msg_to_check_it_0_cnu_14_in_5, msg_to_check_it_0_cnu_42_in_5, msg_to_check_it_0_cnu_70_in_5);
vnu_1 variable_node_167_0(data_167, msg_to_check_it_0_cnu_15_in_5, msg_to_check_it_0_cnu_43_in_5, msg_to_check_it_0_cnu_71_in_5);
vnu_1 variable_node_168_0(data_168, msg_to_check_it_0_cnu_16_in_5, msg_to_check_it_0_cnu_44_in_5, msg_to_check_it_0_cnu_72_in_5);
vnu_1 variable_node_169_0(data_169, msg_to_check_it_0_cnu_17_in_5, msg_to_check_it_0_cnu_45_in_5, msg_to_check_it_0_cnu_73_in_5);
vnu_1 variable_node_170_0(data_170, msg_to_check_it_0_cnu_18_in_5, msg_to_check_it_0_cnu_46_in_5, msg_to_check_it_0_cnu_74_in_5);
vnu_1 variable_node_171_0(data_171, msg_to_check_it_0_cnu_19_in_5, msg_to_check_it_0_cnu_47_in_5, msg_to_check_it_0_cnu_75_in_5);
vnu_1 variable_node_172_0(data_172, msg_to_check_it_0_cnu_20_in_5, msg_to_check_it_0_cnu_48_in_5, msg_to_check_it_0_cnu_76_in_5);
vnu_1 variable_node_173_0(data_173, msg_to_check_it_0_cnu_21_in_5, msg_to_check_it_0_cnu_49_in_5, msg_to_check_it_0_cnu_77_in_5);
vnu_1 variable_node_174_0(data_174, msg_to_check_it_0_cnu_22_in_5, msg_to_check_it_0_cnu_50_in_5, msg_to_check_it_0_cnu_78_in_5);
vnu_1 variable_node_175_0(data_175, msg_to_check_it_0_cnu_23_in_5, msg_to_check_it_0_cnu_51_in_5, msg_to_check_it_0_cnu_79_in_5);
vnu_1 variable_node_176_0(data_176, msg_to_check_it_0_cnu_24_in_5, msg_to_check_it_0_cnu_52_in_5, msg_to_check_it_0_cnu_80_in_5);
vnu_1 variable_node_177_0(data_177, msg_to_check_it_0_cnu_25_in_5, msg_to_check_it_0_cnu_53_in_5, msg_to_check_it_0_cnu_81_in_5);
vnu_1 variable_node_178_0(data_178, msg_to_check_it_0_cnu_26_in_5, msg_to_check_it_0_cnu_54_in_5, msg_to_check_it_0_cnu_82_in_5);
vnu_1 variable_node_179_0(data_179, msg_to_check_it_0_cnu_27_in_5, msg_to_check_it_0_cnu_55_in_5, msg_to_check_it_0_cnu_83_in_5);
vnu_1 variable_node_180_0(data_180, msg_to_check_it_0_cnu_28_in_5, msg_to_check_it_0_cnu_56_in_5, msg_to_check_it_0_cnu_84_in_5);
vnu_1 variable_node_181_0(data_181, msg_to_check_it_0_cnu_29_in_5, msg_to_check_it_0_cnu_57_in_5, msg_to_check_it_0_cnu_85_in_5);
vnu_1 variable_node_182_0(data_182, msg_to_check_it_0_cnu_30_in_5, msg_to_check_it_0_cnu_58_in_5, msg_to_check_it_0_cnu_86_in_5);
vnu_1 variable_node_183_0(data_183, msg_to_check_it_0_cnu_31_in_5, msg_to_check_it_0_cnu_59_in_5, msg_to_check_it_0_cnu_87_in_5);
vnu_1 variable_node_184_0(data_184, msg_to_check_it_0_cnu_32_in_5, msg_to_check_it_0_cnu_60_in_5, msg_to_check_it_0_cnu_88_in_5);
vnu_1 variable_node_185_0(data_185, msg_to_check_it_0_cnu_0_in_5, msg_to_check_it_0_cnu_61_in_5, msg_to_check_it_0_cnu_89_in_5);
vnu_1 variable_node_186_0(data_186, msg_to_check_it_0_cnu_1_in_5, msg_to_check_it_0_cnu_62_in_5, msg_to_check_it_0_cnu_90_in_5);
vnu_1 variable_node_187_0(data_187, msg_to_check_it_0_cnu_2_in_5, msg_to_check_it_0_cnu_63_in_5, msg_to_check_it_0_cnu_91_in_5);
vnu_1 variable_node_188_0(data_188, msg_to_check_it_0_cnu_3_in_5, msg_to_check_it_0_cnu_64_in_5, msg_to_check_it_0_cnu_92_in_5);
vnu_1 variable_node_189_0(data_189, msg_to_check_it_0_cnu_4_in_5, msg_to_check_it_0_cnu_65_in_5, msg_to_check_it_0_cnu_93_in_5);
vnu_1 variable_node_190_0(data_190, msg_to_check_it_0_cnu_5_in_5, msg_to_check_it_0_cnu_33_in_5, msg_to_check_it_0_cnu_94_in_5);
vnu_1 variable_node_191_0(data_191, msg_to_check_it_0_cnu_6_in_5, msg_to_check_it_0_cnu_34_in_5, msg_to_check_it_0_cnu_95_in_5);
vnu_1 variable_node_192_0(data_192, msg_to_check_it_0_cnu_7_in_5, msg_to_check_it_0_cnu_35_in_5, msg_to_check_it_0_cnu_96_in_5);
vnu_1 variable_node_193_0(data_193, msg_to_check_it_0_cnu_8_in_5, msg_to_check_it_0_cnu_36_in_5, msg_to_check_it_0_cnu_97_in_5);
vnu_1 variable_node_194_0(data_194, msg_to_check_it_0_cnu_9_in_5, msg_to_check_it_0_cnu_37_in_5, msg_to_check_it_0_cnu_98_in_5);
vnu_1 variable_node_195_0(data_195, msg_to_check_it_0_cnu_10_in_5, msg_to_check_it_0_cnu_38_in_5, msg_to_check_it_0_cnu_66_in_5);
vnu_1 variable_node_196_0(data_196, msg_to_check_it_0_cnu_11_in_5, msg_to_check_it_0_cnu_39_in_5, msg_to_check_it_0_cnu_67_in_5);
vnu_1 variable_node_197_0(data_197, msg_to_check_it_0_cnu_12_in_5, msg_to_check_it_0_cnu_40_in_5, msg_to_check_it_0_cnu_68_in_5);



cnu check_node_0_0(msg_to_check_it_0_cnu_0_in_0, msg_to_check_it_0_cnu_0_in_1, msg_to_check_it_0_cnu_0_in_2, msg_to_check_it_0_cnu_0_in_3, msg_to_check_it_0_cnu_0_in_4, msg_to_check_it_0_cnu_0_in_5, msg_to_bit_it_1_vnu_2_in_0, msg_to_bit_it_1_vnu_36_in_0, msg_to_bit_it_1_vnu_73_in_0, msg_to_bit_it_1_vnu_108_in_0, msg_to_bit_it_1_vnu_147_in_0, msg_to_bit_it_1_vnu_185_in_0);
cnu check_node_1_0(msg_to_check_it_0_cnu_1_in_0, msg_to_check_it_0_cnu_1_in_1, msg_to_check_it_0_cnu_1_in_2, msg_to_check_it_0_cnu_1_in_3, msg_to_check_it_0_cnu_1_in_4, msg_to_check_it_0_cnu_1_in_5, msg_to_bit_it_1_vnu_3_in_0, msg_to_bit_it_1_vnu_37_in_0, msg_to_bit_it_1_vnu_74_in_0, msg_to_bit_it_1_vnu_109_in_0, msg_to_bit_it_1_vnu_148_in_0, msg_to_bit_it_1_vnu_186_in_0);
cnu check_node_2_0(msg_to_check_it_0_cnu_2_in_0, msg_to_check_it_0_cnu_2_in_1, msg_to_check_it_0_cnu_2_in_2, msg_to_check_it_0_cnu_2_in_3, msg_to_check_it_0_cnu_2_in_4, msg_to_check_it_0_cnu_2_in_5, msg_to_bit_it_1_vnu_4_in_0, msg_to_bit_it_1_vnu_38_in_0, msg_to_bit_it_1_vnu_75_in_0, msg_to_bit_it_1_vnu_110_in_0, msg_to_bit_it_1_vnu_149_in_0, msg_to_bit_it_1_vnu_187_in_0);
cnu check_node_3_0(msg_to_check_it_0_cnu_3_in_0, msg_to_check_it_0_cnu_3_in_1, msg_to_check_it_0_cnu_3_in_2, msg_to_check_it_0_cnu_3_in_3, msg_to_check_it_0_cnu_3_in_4, msg_to_check_it_0_cnu_3_in_5, msg_to_bit_it_1_vnu_5_in_0, msg_to_bit_it_1_vnu_39_in_0, msg_to_bit_it_1_vnu_76_in_0, msg_to_bit_it_1_vnu_111_in_0, msg_to_bit_it_1_vnu_150_in_0, msg_to_bit_it_1_vnu_188_in_0);
cnu check_node_4_0(msg_to_check_it_0_cnu_4_in_0, msg_to_check_it_0_cnu_4_in_1, msg_to_check_it_0_cnu_4_in_2, msg_to_check_it_0_cnu_4_in_3, msg_to_check_it_0_cnu_4_in_4, msg_to_check_it_0_cnu_4_in_5, msg_to_bit_it_1_vnu_6_in_0, msg_to_bit_it_1_vnu_40_in_0, msg_to_bit_it_1_vnu_77_in_0, msg_to_bit_it_1_vnu_112_in_0, msg_to_bit_it_1_vnu_151_in_0, msg_to_bit_it_1_vnu_189_in_0);
cnu check_node_5_0(msg_to_check_it_0_cnu_5_in_0, msg_to_check_it_0_cnu_5_in_1, msg_to_check_it_0_cnu_5_in_2, msg_to_check_it_0_cnu_5_in_3, msg_to_check_it_0_cnu_5_in_4, msg_to_check_it_0_cnu_5_in_5, msg_to_bit_it_1_vnu_7_in_0, msg_to_bit_it_1_vnu_41_in_0, msg_to_bit_it_1_vnu_78_in_0, msg_to_bit_it_1_vnu_113_in_0, msg_to_bit_it_1_vnu_152_in_0, msg_to_bit_it_1_vnu_190_in_0);
cnu check_node_6_0(msg_to_check_it_0_cnu_6_in_0, msg_to_check_it_0_cnu_6_in_1, msg_to_check_it_0_cnu_6_in_2, msg_to_check_it_0_cnu_6_in_3, msg_to_check_it_0_cnu_6_in_4, msg_to_check_it_0_cnu_6_in_5, msg_to_bit_it_1_vnu_8_in_0, msg_to_bit_it_1_vnu_42_in_0, msg_to_bit_it_1_vnu_79_in_0, msg_to_bit_it_1_vnu_114_in_0, msg_to_bit_it_1_vnu_153_in_0, msg_to_bit_it_1_vnu_191_in_0);
cnu check_node_7_0(msg_to_check_it_0_cnu_7_in_0, msg_to_check_it_0_cnu_7_in_1, msg_to_check_it_0_cnu_7_in_2, msg_to_check_it_0_cnu_7_in_3, msg_to_check_it_0_cnu_7_in_4, msg_to_check_it_0_cnu_7_in_5, msg_to_bit_it_1_vnu_9_in_0, msg_to_bit_it_1_vnu_43_in_0, msg_to_bit_it_1_vnu_80_in_0, msg_to_bit_it_1_vnu_115_in_0, msg_to_bit_it_1_vnu_154_in_0, msg_to_bit_it_1_vnu_192_in_0);
cnu check_node_8_0(msg_to_check_it_0_cnu_8_in_0, msg_to_check_it_0_cnu_8_in_1, msg_to_check_it_0_cnu_8_in_2, msg_to_check_it_0_cnu_8_in_3, msg_to_check_it_0_cnu_8_in_4, msg_to_check_it_0_cnu_8_in_5, msg_to_bit_it_1_vnu_10_in_0, msg_to_bit_it_1_vnu_44_in_0, msg_to_bit_it_1_vnu_81_in_0, msg_to_bit_it_1_vnu_116_in_0, msg_to_bit_it_1_vnu_155_in_0, msg_to_bit_it_1_vnu_193_in_0);
cnu check_node_9_0(msg_to_check_it_0_cnu_9_in_0, msg_to_check_it_0_cnu_9_in_1, msg_to_check_it_0_cnu_9_in_2, msg_to_check_it_0_cnu_9_in_3, msg_to_check_it_0_cnu_9_in_4, msg_to_check_it_0_cnu_9_in_5, msg_to_bit_it_1_vnu_11_in_0, msg_to_bit_it_1_vnu_45_in_0, msg_to_bit_it_1_vnu_82_in_0, msg_to_bit_it_1_vnu_117_in_0, msg_to_bit_it_1_vnu_156_in_0, msg_to_bit_it_1_vnu_194_in_0);
cnu check_node_10_0(msg_to_check_it_0_cnu_10_in_0, msg_to_check_it_0_cnu_10_in_1, msg_to_check_it_0_cnu_10_in_2, msg_to_check_it_0_cnu_10_in_3, msg_to_check_it_0_cnu_10_in_4, msg_to_check_it_0_cnu_10_in_5, msg_to_bit_it_1_vnu_12_in_0, msg_to_bit_it_1_vnu_46_in_0, msg_to_bit_it_1_vnu_83_in_0, msg_to_bit_it_1_vnu_118_in_0, msg_to_bit_it_1_vnu_157_in_0, msg_to_bit_it_1_vnu_195_in_0);
cnu check_node_11_0(msg_to_check_it_0_cnu_11_in_0, msg_to_check_it_0_cnu_11_in_1, msg_to_check_it_0_cnu_11_in_2, msg_to_check_it_0_cnu_11_in_3, msg_to_check_it_0_cnu_11_in_4, msg_to_check_it_0_cnu_11_in_5, msg_to_bit_it_1_vnu_13_in_0, msg_to_bit_it_1_vnu_47_in_0, msg_to_bit_it_1_vnu_84_in_0, msg_to_bit_it_1_vnu_119_in_0, msg_to_bit_it_1_vnu_158_in_0, msg_to_bit_it_1_vnu_196_in_0);
cnu check_node_12_0(msg_to_check_it_0_cnu_12_in_0, msg_to_check_it_0_cnu_12_in_1, msg_to_check_it_0_cnu_12_in_2, msg_to_check_it_0_cnu_12_in_3, msg_to_check_it_0_cnu_12_in_4, msg_to_check_it_0_cnu_12_in_5, msg_to_bit_it_1_vnu_14_in_0, msg_to_bit_it_1_vnu_48_in_0, msg_to_bit_it_1_vnu_85_in_0, msg_to_bit_it_1_vnu_120_in_0, msg_to_bit_it_1_vnu_159_in_0, msg_to_bit_it_1_vnu_197_in_0);
cnu check_node_13_0(msg_to_check_it_0_cnu_13_in_0, msg_to_check_it_0_cnu_13_in_1, msg_to_check_it_0_cnu_13_in_2, msg_to_check_it_0_cnu_13_in_3, msg_to_check_it_0_cnu_13_in_4, msg_to_check_it_0_cnu_13_in_5, msg_to_bit_it_1_vnu_15_in_0, msg_to_bit_it_1_vnu_49_in_0, msg_to_bit_it_1_vnu_86_in_0, msg_to_bit_it_1_vnu_121_in_0, msg_to_bit_it_1_vnu_160_in_0, msg_to_bit_it_1_vnu_165_in_0);
cnu check_node_14_0(msg_to_check_it_0_cnu_14_in_0, msg_to_check_it_0_cnu_14_in_1, msg_to_check_it_0_cnu_14_in_2, msg_to_check_it_0_cnu_14_in_3, msg_to_check_it_0_cnu_14_in_4, msg_to_check_it_0_cnu_14_in_5, msg_to_bit_it_1_vnu_16_in_0, msg_to_bit_it_1_vnu_50_in_0, msg_to_bit_it_1_vnu_87_in_0, msg_to_bit_it_1_vnu_122_in_0, msg_to_bit_it_1_vnu_161_in_0, msg_to_bit_it_1_vnu_166_in_0);
cnu check_node_15_0(msg_to_check_it_0_cnu_15_in_0, msg_to_check_it_0_cnu_15_in_1, msg_to_check_it_0_cnu_15_in_2, msg_to_check_it_0_cnu_15_in_3, msg_to_check_it_0_cnu_15_in_4, msg_to_check_it_0_cnu_15_in_5, msg_to_bit_it_1_vnu_17_in_0, msg_to_bit_it_1_vnu_51_in_0, msg_to_bit_it_1_vnu_88_in_0, msg_to_bit_it_1_vnu_123_in_0, msg_to_bit_it_1_vnu_162_in_0, msg_to_bit_it_1_vnu_167_in_0);
cnu check_node_16_0(msg_to_check_it_0_cnu_16_in_0, msg_to_check_it_0_cnu_16_in_1, msg_to_check_it_0_cnu_16_in_2, msg_to_check_it_0_cnu_16_in_3, msg_to_check_it_0_cnu_16_in_4, msg_to_check_it_0_cnu_16_in_5, msg_to_bit_it_1_vnu_18_in_0, msg_to_bit_it_1_vnu_52_in_0, msg_to_bit_it_1_vnu_89_in_0, msg_to_bit_it_1_vnu_124_in_0, msg_to_bit_it_1_vnu_163_in_0, msg_to_bit_it_1_vnu_168_in_0);
cnu check_node_17_0(msg_to_check_it_0_cnu_17_in_0, msg_to_check_it_0_cnu_17_in_1, msg_to_check_it_0_cnu_17_in_2, msg_to_check_it_0_cnu_17_in_3, msg_to_check_it_0_cnu_17_in_4, msg_to_check_it_0_cnu_17_in_5, msg_to_bit_it_1_vnu_19_in_0, msg_to_bit_it_1_vnu_53_in_0, msg_to_bit_it_1_vnu_90_in_0, msg_to_bit_it_1_vnu_125_in_0, msg_to_bit_it_1_vnu_164_in_0, msg_to_bit_it_1_vnu_169_in_0);
cnu check_node_18_0(msg_to_check_it_0_cnu_18_in_0, msg_to_check_it_0_cnu_18_in_1, msg_to_check_it_0_cnu_18_in_2, msg_to_check_it_0_cnu_18_in_3, msg_to_check_it_0_cnu_18_in_4, msg_to_check_it_0_cnu_18_in_5, msg_to_bit_it_1_vnu_20_in_0, msg_to_bit_it_1_vnu_54_in_0, msg_to_bit_it_1_vnu_91_in_0, msg_to_bit_it_1_vnu_126_in_0, msg_to_bit_it_1_vnu_132_in_0, msg_to_bit_it_1_vnu_170_in_0);
cnu check_node_19_0(msg_to_check_it_0_cnu_19_in_0, msg_to_check_it_0_cnu_19_in_1, msg_to_check_it_0_cnu_19_in_2, msg_to_check_it_0_cnu_19_in_3, msg_to_check_it_0_cnu_19_in_4, msg_to_check_it_0_cnu_19_in_5, msg_to_bit_it_1_vnu_21_in_0, msg_to_bit_it_1_vnu_55_in_0, msg_to_bit_it_1_vnu_92_in_0, msg_to_bit_it_1_vnu_127_in_0, msg_to_bit_it_1_vnu_133_in_0, msg_to_bit_it_1_vnu_171_in_0);
cnu check_node_20_0(msg_to_check_it_0_cnu_20_in_0, msg_to_check_it_0_cnu_20_in_1, msg_to_check_it_0_cnu_20_in_2, msg_to_check_it_0_cnu_20_in_3, msg_to_check_it_0_cnu_20_in_4, msg_to_check_it_0_cnu_20_in_5, msg_to_bit_it_1_vnu_22_in_0, msg_to_bit_it_1_vnu_56_in_0, msg_to_bit_it_1_vnu_93_in_0, msg_to_bit_it_1_vnu_128_in_0, msg_to_bit_it_1_vnu_134_in_0, msg_to_bit_it_1_vnu_172_in_0);
cnu check_node_21_0(msg_to_check_it_0_cnu_21_in_0, msg_to_check_it_0_cnu_21_in_1, msg_to_check_it_0_cnu_21_in_2, msg_to_check_it_0_cnu_21_in_3, msg_to_check_it_0_cnu_21_in_4, msg_to_check_it_0_cnu_21_in_5, msg_to_bit_it_1_vnu_23_in_0, msg_to_bit_it_1_vnu_57_in_0, msg_to_bit_it_1_vnu_94_in_0, msg_to_bit_it_1_vnu_129_in_0, msg_to_bit_it_1_vnu_135_in_0, msg_to_bit_it_1_vnu_173_in_0);
cnu check_node_22_0(msg_to_check_it_0_cnu_22_in_0, msg_to_check_it_0_cnu_22_in_1, msg_to_check_it_0_cnu_22_in_2, msg_to_check_it_0_cnu_22_in_3, msg_to_check_it_0_cnu_22_in_4, msg_to_check_it_0_cnu_22_in_5, msg_to_bit_it_1_vnu_24_in_0, msg_to_bit_it_1_vnu_58_in_0, msg_to_bit_it_1_vnu_95_in_0, msg_to_bit_it_1_vnu_130_in_0, msg_to_bit_it_1_vnu_136_in_0, msg_to_bit_it_1_vnu_174_in_0);
cnu check_node_23_0(msg_to_check_it_0_cnu_23_in_0, msg_to_check_it_0_cnu_23_in_1, msg_to_check_it_0_cnu_23_in_2, msg_to_check_it_0_cnu_23_in_3, msg_to_check_it_0_cnu_23_in_4, msg_to_check_it_0_cnu_23_in_5, msg_to_bit_it_1_vnu_25_in_0, msg_to_bit_it_1_vnu_59_in_0, msg_to_bit_it_1_vnu_96_in_0, msg_to_bit_it_1_vnu_131_in_0, msg_to_bit_it_1_vnu_137_in_0, msg_to_bit_it_1_vnu_175_in_0);
cnu check_node_24_0(msg_to_check_it_0_cnu_24_in_0, msg_to_check_it_0_cnu_24_in_1, msg_to_check_it_0_cnu_24_in_2, msg_to_check_it_0_cnu_24_in_3, msg_to_check_it_0_cnu_24_in_4, msg_to_check_it_0_cnu_24_in_5, msg_to_bit_it_1_vnu_26_in_0, msg_to_bit_it_1_vnu_60_in_0, msg_to_bit_it_1_vnu_97_in_0, msg_to_bit_it_1_vnu_99_in_0, msg_to_bit_it_1_vnu_138_in_0, msg_to_bit_it_1_vnu_176_in_0);
cnu check_node_25_0(msg_to_check_it_0_cnu_25_in_0, msg_to_check_it_0_cnu_25_in_1, msg_to_check_it_0_cnu_25_in_2, msg_to_check_it_0_cnu_25_in_3, msg_to_check_it_0_cnu_25_in_4, msg_to_check_it_0_cnu_25_in_5, msg_to_bit_it_1_vnu_27_in_0, msg_to_bit_it_1_vnu_61_in_0, msg_to_bit_it_1_vnu_98_in_0, msg_to_bit_it_1_vnu_100_in_0, msg_to_bit_it_1_vnu_139_in_0, msg_to_bit_it_1_vnu_177_in_0);
cnu check_node_26_0(msg_to_check_it_0_cnu_26_in_0, msg_to_check_it_0_cnu_26_in_1, msg_to_check_it_0_cnu_26_in_2, msg_to_check_it_0_cnu_26_in_3, msg_to_check_it_0_cnu_26_in_4, msg_to_check_it_0_cnu_26_in_5, msg_to_bit_it_1_vnu_28_in_0, msg_to_bit_it_1_vnu_62_in_0, msg_to_bit_it_1_vnu_66_in_0, msg_to_bit_it_1_vnu_101_in_0, msg_to_bit_it_1_vnu_140_in_0, msg_to_bit_it_1_vnu_178_in_0);
cnu check_node_27_0(msg_to_check_it_0_cnu_27_in_0, msg_to_check_it_0_cnu_27_in_1, msg_to_check_it_0_cnu_27_in_2, msg_to_check_it_0_cnu_27_in_3, msg_to_check_it_0_cnu_27_in_4, msg_to_check_it_0_cnu_27_in_5, msg_to_bit_it_1_vnu_29_in_0, msg_to_bit_it_1_vnu_63_in_0, msg_to_bit_it_1_vnu_67_in_0, msg_to_bit_it_1_vnu_102_in_0, msg_to_bit_it_1_vnu_141_in_0, msg_to_bit_it_1_vnu_179_in_0);
cnu check_node_28_0(msg_to_check_it_0_cnu_28_in_0, msg_to_check_it_0_cnu_28_in_1, msg_to_check_it_0_cnu_28_in_2, msg_to_check_it_0_cnu_28_in_3, msg_to_check_it_0_cnu_28_in_4, msg_to_check_it_0_cnu_28_in_5, msg_to_bit_it_1_vnu_30_in_0, msg_to_bit_it_1_vnu_64_in_0, msg_to_bit_it_1_vnu_68_in_0, msg_to_bit_it_1_vnu_103_in_0, msg_to_bit_it_1_vnu_142_in_0, msg_to_bit_it_1_vnu_180_in_0);
cnu check_node_29_0(msg_to_check_it_0_cnu_29_in_0, msg_to_check_it_0_cnu_29_in_1, msg_to_check_it_0_cnu_29_in_2, msg_to_check_it_0_cnu_29_in_3, msg_to_check_it_0_cnu_29_in_4, msg_to_check_it_0_cnu_29_in_5, msg_to_bit_it_1_vnu_31_in_0, msg_to_bit_it_1_vnu_65_in_0, msg_to_bit_it_1_vnu_69_in_0, msg_to_bit_it_1_vnu_104_in_0, msg_to_bit_it_1_vnu_143_in_0, msg_to_bit_it_1_vnu_181_in_0);
cnu check_node_30_0(msg_to_check_it_0_cnu_30_in_0, msg_to_check_it_0_cnu_30_in_1, msg_to_check_it_0_cnu_30_in_2, msg_to_check_it_0_cnu_30_in_3, msg_to_check_it_0_cnu_30_in_4, msg_to_check_it_0_cnu_30_in_5, msg_to_bit_it_1_vnu_32_in_0, msg_to_bit_it_1_vnu_33_in_0, msg_to_bit_it_1_vnu_70_in_0, msg_to_bit_it_1_vnu_105_in_0, msg_to_bit_it_1_vnu_144_in_0, msg_to_bit_it_1_vnu_182_in_0);
cnu check_node_31_0(msg_to_check_it_0_cnu_31_in_0, msg_to_check_it_0_cnu_31_in_1, msg_to_check_it_0_cnu_31_in_2, msg_to_check_it_0_cnu_31_in_3, msg_to_check_it_0_cnu_31_in_4, msg_to_check_it_0_cnu_31_in_5, msg_to_bit_it_1_vnu_0_in_0, msg_to_bit_it_1_vnu_34_in_0, msg_to_bit_it_1_vnu_71_in_0, msg_to_bit_it_1_vnu_106_in_0, msg_to_bit_it_1_vnu_145_in_0, msg_to_bit_it_1_vnu_183_in_0);
cnu check_node_32_0(msg_to_check_it_0_cnu_32_in_0, msg_to_check_it_0_cnu_32_in_1, msg_to_check_it_0_cnu_32_in_2, msg_to_check_it_0_cnu_32_in_3, msg_to_check_it_0_cnu_32_in_4, msg_to_check_it_0_cnu_32_in_5, msg_to_bit_it_1_vnu_1_in_0, msg_to_bit_it_1_vnu_35_in_0, msg_to_bit_it_1_vnu_72_in_0, msg_to_bit_it_1_vnu_107_in_0, msg_to_bit_it_1_vnu_146_in_0, msg_to_bit_it_1_vnu_184_in_0);
cnu check_node_33_0(msg_to_check_it_0_cnu_33_in_0, msg_to_check_it_0_cnu_33_in_1, msg_to_check_it_0_cnu_33_in_2, msg_to_check_it_0_cnu_33_in_3, msg_to_check_it_0_cnu_33_in_4, msg_to_check_it_0_cnu_33_in_5, msg_to_bit_it_1_vnu_4_in_1, msg_to_bit_it_1_vnu_38_in_1, msg_to_bit_it_1_vnu_77_in_1, msg_to_bit_it_1_vnu_111_in_1, msg_to_bit_it_1_vnu_155_in_1, msg_to_bit_it_1_vnu_190_in_1);
cnu check_node_34_0(msg_to_check_it_0_cnu_34_in_0, msg_to_check_it_0_cnu_34_in_1, msg_to_check_it_0_cnu_34_in_2, msg_to_check_it_0_cnu_34_in_3, msg_to_check_it_0_cnu_34_in_4, msg_to_check_it_0_cnu_34_in_5, msg_to_bit_it_1_vnu_5_in_1, msg_to_bit_it_1_vnu_39_in_1, msg_to_bit_it_1_vnu_78_in_1, msg_to_bit_it_1_vnu_112_in_1, msg_to_bit_it_1_vnu_156_in_1, msg_to_bit_it_1_vnu_191_in_1);
cnu check_node_35_0(msg_to_check_it_0_cnu_35_in_0, msg_to_check_it_0_cnu_35_in_1, msg_to_check_it_0_cnu_35_in_2, msg_to_check_it_0_cnu_35_in_3, msg_to_check_it_0_cnu_35_in_4, msg_to_check_it_0_cnu_35_in_5, msg_to_bit_it_1_vnu_6_in_1, msg_to_bit_it_1_vnu_40_in_1, msg_to_bit_it_1_vnu_79_in_1, msg_to_bit_it_1_vnu_113_in_1, msg_to_bit_it_1_vnu_157_in_1, msg_to_bit_it_1_vnu_192_in_1);
cnu check_node_36_0(msg_to_check_it_0_cnu_36_in_0, msg_to_check_it_0_cnu_36_in_1, msg_to_check_it_0_cnu_36_in_2, msg_to_check_it_0_cnu_36_in_3, msg_to_check_it_0_cnu_36_in_4, msg_to_check_it_0_cnu_36_in_5, msg_to_bit_it_1_vnu_7_in_1, msg_to_bit_it_1_vnu_41_in_1, msg_to_bit_it_1_vnu_80_in_1, msg_to_bit_it_1_vnu_114_in_1, msg_to_bit_it_1_vnu_158_in_1, msg_to_bit_it_1_vnu_193_in_1);
cnu check_node_37_0(msg_to_check_it_0_cnu_37_in_0, msg_to_check_it_0_cnu_37_in_1, msg_to_check_it_0_cnu_37_in_2, msg_to_check_it_0_cnu_37_in_3, msg_to_check_it_0_cnu_37_in_4, msg_to_check_it_0_cnu_37_in_5, msg_to_bit_it_1_vnu_8_in_1, msg_to_bit_it_1_vnu_42_in_1, msg_to_bit_it_1_vnu_81_in_1, msg_to_bit_it_1_vnu_115_in_1, msg_to_bit_it_1_vnu_159_in_1, msg_to_bit_it_1_vnu_194_in_1);
cnu check_node_38_0(msg_to_check_it_0_cnu_38_in_0, msg_to_check_it_0_cnu_38_in_1, msg_to_check_it_0_cnu_38_in_2, msg_to_check_it_0_cnu_38_in_3, msg_to_check_it_0_cnu_38_in_4, msg_to_check_it_0_cnu_38_in_5, msg_to_bit_it_1_vnu_9_in_1, msg_to_bit_it_1_vnu_43_in_1, msg_to_bit_it_1_vnu_82_in_1, msg_to_bit_it_1_vnu_116_in_1, msg_to_bit_it_1_vnu_160_in_1, msg_to_bit_it_1_vnu_195_in_1);
cnu check_node_39_0(msg_to_check_it_0_cnu_39_in_0, msg_to_check_it_0_cnu_39_in_1, msg_to_check_it_0_cnu_39_in_2, msg_to_check_it_0_cnu_39_in_3, msg_to_check_it_0_cnu_39_in_4, msg_to_check_it_0_cnu_39_in_5, msg_to_bit_it_1_vnu_10_in_1, msg_to_bit_it_1_vnu_44_in_1, msg_to_bit_it_1_vnu_83_in_1, msg_to_bit_it_1_vnu_117_in_1, msg_to_bit_it_1_vnu_161_in_1, msg_to_bit_it_1_vnu_196_in_1);
cnu check_node_40_0(msg_to_check_it_0_cnu_40_in_0, msg_to_check_it_0_cnu_40_in_1, msg_to_check_it_0_cnu_40_in_2, msg_to_check_it_0_cnu_40_in_3, msg_to_check_it_0_cnu_40_in_4, msg_to_check_it_0_cnu_40_in_5, msg_to_bit_it_1_vnu_11_in_1, msg_to_bit_it_1_vnu_45_in_1, msg_to_bit_it_1_vnu_84_in_1, msg_to_bit_it_1_vnu_118_in_1, msg_to_bit_it_1_vnu_162_in_1, msg_to_bit_it_1_vnu_197_in_1);
cnu check_node_41_0(msg_to_check_it_0_cnu_41_in_0, msg_to_check_it_0_cnu_41_in_1, msg_to_check_it_0_cnu_41_in_2, msg_to_check_it_0_cnu_41_in_3, msg_to_check_it_0_cnu_41_in_4, msg_to_check_it_0_cnu_41_in_5, msg_to_bit_it_1_vnu_12_in_1, msg_to_bit_it_1_vnu_46_in_1, msg_to_bit_it_1_vnu_85_in_1, msg_to_bit_it_1_vnu_119_in_1, msg_to_bit_it_1_vnu_163_in_1, msg_to_bit_it_1_vnu_165_in_1);
cnu check_node_42_0(msg_to_check_it_0_cnu_42_in_0, msg_to_check_it_0_cnu_42_in_1, msg_to_check_it_0_cnu_42_in_2, msg_to_check_it_0_cnu_42_in_3, msg_to_check_it_0_cnu_42_in_4, msg_to_check_it_0_cnu_42_in_5, msg_to_bit_it_1_vnu_13_in_1, msg_to_bit_it_1_vnu_47_in_1, msg_to_bit_it_1_vnu_86_in_1, msg_to_bit_it_1_vnu_120_in_1, msg_to_bit_it_1_vnu_164_in_1, msg_to_bit_it_1_vnu_166_in_1);
cnu check_node_43_0(msg_to_check_it_0_cnu_43_in_0, msg_to_check_it_0_cnu_43_in_1, msg_to_check_it_0_cnu_43_in_2, msg_to_check_it_0_cnu_43_in_3, msg_to_check_it_0_cnu_43_in_4, msg_to_check_it_0_cnu_43_in_5, msg_to_bit_it_1_vnu_14_in_1, msg_to_bit_it_1_vnu_48_in_1, msg_to_bit_it_1_vnu_87_in_1, msg_to_bit_it_1_vnu_121_in_1, msg_to_bit_it_1_vnu_132_in_1, msg_to_bit_it_1_vnu_167_in_1);
cnu check_node_44_0(msg_to_check_it_0_cnu_44_in_0, msg_to_check_it_0_cnu_44_in_1, msg_to_check_it_0_cnu_44_in_2, msg_to_check_it_0_cnu_44_in_3, msg_to_check_it_0_cnu_44_in_4, msg_to_check_it_0_cnu_44_in_5, msg_to_bit_it_1_vnu_15_in_1, msg_to_bit_it_1_vnu_49_in_1, msg_to_bit_it_1_vnu_88_in_1, msg_to_bit_it_1_vnu_122_in_1, msg_to_bit_it_1_vnu_133_in_1, msg_to_bit_it_1_vnu_168_in_1);
cnu check_node_45_0(msg_to_check_it_0_cnu_45_in_0, msg_to_check_it_0_cnu_45_in_1, msg_to_check_it_0_cnu_45_in_2, msg_to_check_it_0_cnu_45_in_3, msg_to_check_it_0_cnu_45_in_4, msg_to_check_it_0_cnu_45_in_5, msg_to_bit_it_1_vnu_16_in_1, msg_to_bit_it_1_vnu_50_in_1, msg_to_bit_it_1_vnu_89_in_1, msg_to_bit_it_1_vnu_123_in_1, msg_to_bit_it_1_vnu_134_in_1, msg_to_bit_it_1_vnu_169_in_1);
cnu check_node_46_0(msg_to_check_it_0_cnu_46_in_0, msg_to_check_it_0_cnu_46_in_1, msg_to_check_it_0_cnu_46_in_2, msg_to_check_it_0_cnu_46_in_3, msg_to_check_it_0_cnu_46_in_4, msg_to_check_it_0_cnu_46_in_5, msg_to_bit_it_1_vnu_17_in_1, msg_to_bit_it_1_vnu_51_in_1, msg_to_bit_it_1_vnu_90_in_1, msg_to_bit_it_1_vnu_124_in_1, msg_to_bit_it_1_vnu_135_in_1, msg_to_bit_it_1_vnu_170_in_1);
cnu check_node_47_0(msg_to_check_it_0_cnu_47_in_0, msg_to_check_it_0_cnu_47_in_1, msg_to_check_it_0_cnu_47_in_2, msg_to_check_it_0_cnu_47_in_3, msg_to_check_it_0_cnu_47_in_4, msg_to_check_it_0_cnu_47_in_5, msg_to_bit_it_1_vnu_18_in_1, msg_to_bit_it_1_vnu_52_in_1, msg_to_bit_it_1_vnu_91_in_1, msg_to_bit_it_1_vnu_125_in_1, msg_to_bit_it_1_vnu_136_in_1, msg_to_bit_it_1_vnu_171_in_1);
cnu check_node_48_0(msg_to_check_it_0_cnu_48_in_0, msg_to_check_it_0_cnu_48_in_1, msg_to_check_it_0_cnu_48_in_2, msg_to_check_it_0_cnu_48_in_3, msg_to_check_it_0_cnu_48_in_4, msg_to_check_it_0_cnu_48_in_5, msg_to_bit_it_1_vnu_19_in_1, msg_to_bit_it_1_vnu_53_in_1, msg_to_bit_it_1_vnu_92_in_1, msg_to_bit_it_1_vnu_126_in_1, msg_to_bit_it_1_vnu_137_in_1, msg_to_bit_it_1_vnu_172_in_1);
cnu check_node_49_0(msg_to_check_it_0_cnu_49_in_0, msg_to_check_it_0_cnu_49_in_1, msg_to_check_it_0_cnu_49_in_2, msg_to_check_it_0_cnu_49_in_3, msg_to_check_it_0_cnu_49_in_4, msg_to_check_it_0_cnu_49_in_5, msg_to_bit_it_1_vnu_20_in_1, msg_to_bit_it_1_vnu_54_in_1, msg_to_bit_it_1_vnu_93_in_1, msg_to_bit_it_1_vnu_127_in_1, msg_to_bit_it_1_vnu_138_in_1, msg_to_bit_it_1_vnu_173_in_1);
cnu check_node_50_0(msg_to_check_it_0_cnu_50_in_0, msg_to_check_it_0_cnu_50_in_1, msg_to_check_it_0_cnu_50_in_2, msg_to_check_it_0_cnu_50_in_3, msg_to_check_it_0_cnu_50_in_4, msg_to_check_it_0_cnu_50_in_5, msg_to_bit_it_1_vnu_21_in_1, msg_to_bit_it_1_vnu_55_in_1, msg_to_bit_it_1_vnu_94_in_1, msg_to_bit_it_1_vnu_128_in_1, msg_to_bit_it_1_vnu_139_in_1, msg_to_bit_it_1_vnu_174_in_1);
cnu check_node_51_0(msg_to_check_it_0_cnu_51_in_0, msg_to_check_it_0_cnu_51_in_1, msg_to_check_it_0_cnu_51_in_2, msg_to_check_it_0_cnu_51_in_3, msg_to_check_it_0_cnu_51_in_4, msg_to_check_it_0_cnu_51_in_5, msg_to_bit_it_1_vnu_22_in_1, msg_to_bit_it_1_vnu_56_in_1, msg_to_bit_it_1_vnu_95_in_1, msg_to_bit_it_1_vnu_129_in_1, msg_to_bit_it_1_vnu_140_in_1, msg_to_bit_it_1_vnu_175_in_1);
cnu check_node_52_0(msg_to_check_it_0_cnu_52_in_0, msg_to_check_it_0_cnu_52_in_1, msg_to_check_it_0_cnu_52_in_2, msg_to_check_it_0_cnu_52_in_3, msg_to_check_it_0_cnu_52_in_4, msg_to_check_it_0_cnu_52_in_5, msg_to_bit_it_1_vnu_23_in_1, msg_to_bit_it_1_vnu_57_in_1, msg_to_bit_it_1_vnu_96_in_1, msg_to_bit_it_1_vnu_130_in_1, msg_to_bit_it_1_vnu_141_in_1, msg_to_bit_it_1_vnu_176_in_1);
cnu check_node_53_0(msg_to_check_it_0_cnu_53_in_0, msg_to_check_it_0_cnu_53_in_1, msg_to_check_it_0_cnu_53_in_2, msg_to_check_it_0_cnu_53_in_3, msg_to_check_it_0_cnu_53_in_4, msg_to_check_it_0_cnu_53_in_5, msg_to_bit_it_1_vnu_24_in_1, msg_to_bit_it_1_vnu_58_in_1, msg_to_bit_it_1_vnu_97_in_1, msg_to_bit_it_1_vnu_131_in_1, msg_to_bit_it_1_vnu_142_in_1, msg_to_bit_it_1_vnu_177_in_1);
cnu check_node_54_0(msg_to_check_it_0_cnu_54_in_0, msg_to_check_it_0_cnu_54_in_1, msg_to_check_it_0_cnu_54_in_2, msg_to_check_it_0_cnu_54_in_3, msg_to_check_it_0_cnu_54_in_4, msg_to_check_it_0_cnu_54_in_5, msg_to_bit_it_1_vnu_25_in_1, msg_to_bit_it_1_vnu_59_in_1, msg_to_bit_it_1_vnu_98_in_1, msg_to_bit_it_1_vnu_99_in_1, msg_to_bit_it_1_vnu_143_in_1, msg_to_bit_it_1_vnu_178_in_1);
cnu check_node_55_0(msg_to_check_it_0_cnu_55_in_0, msg_to_check_it_0_cnu_55_in_1, msg_to_check_it_0_cnu_55_in_2, msg_to_check_it_0_cnu_55_in_3, msg_to_check_it_0_cnu_55_in_4, msg_to_check_it_0_cnu_55_in_5, msg_to_bit_it_1_vnu_26_in_1, msg_to_bit_it_1_vnu_60_in_1, msg_to_bit_it_1_vnu_66_in_1, msg_to_bit_it_1_vnu_100_in_1, msg_to_bit_it_1_vnu_144_in_1, msg_to_bit_it_1_vnu_179_in_1);
cnu check_node_56_0(msg_to_check_it_0_cnu_56_in_0, msg_to_check_it_0_cnu_56_in_1, msg_to_check_it_0_cnu_56_in_2, msg_to_check_it_0_cnu_56_in_3, msg_to_check_it_0_cnu_56_in_4, msg_to_check_it_0_cnu_56_in_5, msg_to_bit_it_1_vnu_27_in_1, msg_to_bit_it_1_vnu_61_in_1, msg_to_bit_it_1_vnu_67_in_1, msg_to_bit_it_1_vnu_101_in_1, msg_to_bit_it_1_vnu_145_in_1, msg_to_bit_it_1_vnu_180_in_1);
cnu check_node_57_0(msg_to_check_it_0_cnu_57_in_0, msg_to_check_it_0_cnu_57_in_1, msg_to_check_it_0_cnu_57_in_2, msg_to_check_it_0_cnu_57_in_3, msg_to_check_it_0_cnu_57_in_4, msg_to_check_it_0_cnu_57_in_5, msg_to_bit_it_1_vnu_28_in_1, msg_to_bit_it_1_vnu_62_in_1, msg_to_bit_it_1_vnu_68_in_1, msg_to_bit_it_1_vnu_102_in_1, msg_to_bit_it_1_vnu_146_in_1, msg_to_bit_it_1_vnu_181_in_1);
cnu check_node_58_0(msg_to_check_it_0_cnu_58_in_0, msg_to_check_it_0_cnu_58_in_1, msg_to_check_it_0_cnu_58_in_2, msg_to_check_it_0_cnu_58_in_3, msg_to_check_it_0_cnu_58_in_4, msg_to_check_it_0_cnu_58_in_5, msg_to_bit_it_1_vnu_29_in_1, msg_to_bit_it_1_vnu_63_in_1, msg_to_bit_it_1_vnu_69_in_1, msg_to_bit_it_1_vnu_103_in_1, msg_to_bit_it_1_vnu_147_in_1, msg_to_bit_it_1_vnu_182_in_1);
cnu check_node_59_0(msg_to_check_it_0_cnu_59_in_0, msg_to_check_it_0_cnu_59_in_1, msg_to_check_it_0_cnu_59_in_2, msg_to_check_it_0_cnu_59_in_3, msg_to_check_it_0_cnu_59_in_4, msg_to_check_it_0_cnu_59_in_5, msg_to_bit_it_1_vnu_30_in_1, msg_to_bit_it_1_vnu_64_in_1, msg_to_bit_it_1_vnu_70_in_1, msg_to_bit_it_1_vnu_104_in_1, msg_to_bit_it_1_vnu_148_in_1, msg_to_bit_it_1_vnu_183_in_1);
cnu check_node_60_0(msg_to_check_it_0_cnu_60_in_0, msg_to_check_it_0_cnu_60_in_1, msg_to_check_it_0_cnu_60_in_2, msg_to_check_it_0_cnu_60_in_3, msg_to_check_it_0_cnu_60_in_4, msg_to_check_it_0_cnu_60_in_5, msg_to_bit_it_1_vnu_31_in_1, msg_to_bit_it_1_vnu_65_in_1, msg_to_bit_it_1_vnu_71_in_1, msg_to_bit_it_1_vnu_105_in_1, msg_to_bit_it_1_vnu_149_in_1, msg_to_bit_it_1_vnu_184_in_1);
cnu check_node_61_0(msg_to_check_it_0_cnu_61_in_0, msg_to_check_it_0_cnu_61_in_1, msg_to_check_it_0_cnu_61_in_2, msg_to_check_it_0_cnu_61_in_3, msg_to_check_it_0_cnu_61_in_4, msg_to_check_it_0_cnu_61_in_5, msg_to_bit_it_1_vnu_32_in_1, msg_to_bit_it_1_vnu_33_in_1, msg_to_bit_it_1_vnu_72_in_1, msg_to_bit_it_1_vnu_106_in_1, msg_to_bit_it_1_vnu_150_in_1, msg_to_bit_it_1_vnu_185_in_1);
cnu check_node_62_0(msg_to_check_it_0_cnu_62_in_0, msg_to_check_it_0_cnu_62_in_1, msg_to_check_it_0_cnu_62_in_2, msg_to_check_it_0_cnu_62_in_3, msg_to_check_it_0_cnu_62_in_4, msg_to_check_it_0_cnu_62_in_5, msg_to_bit_it_1_vnu_0_in_1, msg_to_bit_it_1_vnu_34_in_1, msg_to_bit_it_1_vnu_73_in_1, msg_to_bit_it_1_vnu_107_in_1, msg_to_bit_it_1_vnu_151_in_1, msg_to_bit_it_1_vnu_186_in_1);
cnu check_node_63_0(msg_to_check_it_0_cnu_63_in_0, msg_to_check_it_0_cnu_63_in_1, msg_to_check_it_0_cnu_63_in_2, msg_to_check_it_0_cnu_63_in_3, msg_to_check_it_0_cnu_63_in_4, msg_to_check_it_0_cnu_63_in_5, msg_to_bit_it_1_vnu_1_in_1, msg_to_bit_it_1_vnu_35_in_1, msg_to_bit_it_1_vnu_74_in_1, msg_to_bit_it_1_vnu_108_in_1, msg_to_bit_it_1_vnu_152_in_1, msg_to_bit_it_1_vnu_187_in_1);
cnu check_node_64_0(msg_to_check_it_0_cnu_64_in_0, msg_to_check_it_0_cnu_64_in_1, msg_to_check_it_0_cnu_64_in_2, msg_to_check_it_0_cnu_64_in_3, msg_to_check_it_0_cnu_64_in_4, msg_to_check_it_0_cnu_64_in_5, msg_to_bit_it_1_vnu_2_in_1, msg_to_bit_it_1_vnu_36_in_1, msg_to_bit_it_1_vnu_75_in_1, msg_to_bit_it_1_vnu_109_in_1, msg_to_bit_it_1_vnu_153_in_1, msg_to_bit_it_1_vnu_188_in_1);
cnu check_node_65_0(msg_to_check_it_0_cnu_65_in_0, msg_to_check_it_0_cnu_65_in_1, msg_to_check_it_0_cnu_65_in_2, msg_to_check_it_0_cnu_65_in_3, msg_to_check_it_0_cnu_65_in_4, msg_to_check_it_0_cnu_65_in_5, msg_to_bit_it_1_vnu_3_in_1, msg_to_bit_it_1_vnu_37_in_1, msg_to_bit_it_1_vnu_76_in_1, msg_to_bit_it_1_vnu_110_in_1, msg_to_bit_it_1_vnu_154_in_1, msg_to_bit_it_1_vnu_189_in_1);
cnu check_node_66_0(msg_to_check_it_0_cnu_66_in_0, msg_to_check_it_0_cnu_66_in_1, msg_to_check_it_0_cnu_66_in_2, msg_to_check_it_0_cnu_66_in_3, msg_to_check_it_0_cnu_66_in_4, msg_to_check_it_0_cnu_66_in_5, msg_to_bit_it_1_vnu_6_in_2, msg_to_bit_it_1_vnu_41_in_2, msg_to_bit_it_1_vnu_80_in_2, msg_to_bit_it_1_vnu_118_in_2, msg_to_bit_it_1_vnu_159_in_2, msg_to_bit_it_1_vnu_195_in_2);
cnu check_node_67_0(msg_to_check_it_0_cnu_67_in_0, msg_to_check_it_0_cnu_67_in_1, msg_to_check_it_0_cnu_67_in_2, msg_to_check_it_0_cnu_67_in_3, msg_to_check_it_0_cnu_67_in_4, msg_to_check_it_0_cnu_67_in_5, msg_to_bit_it_1_vnu_7_in_2, msg_to_bit_it_1_vnu_42_in_2, msg_to_bit_it_1_vnu_81_in_2, msg_to_bit_it_1_vnu_119_in_2, msg_to_bit_it_1_vnu_160_in_2, msg_to_bit_it_1_vnu_196_in_2);
cnu check_node_68_0(msg_to_check_it_0_cnu_68_in_0, msg_to_check_it_0_cnu_68_in_1, msg_to_check_it_0_cnu_68_in_2, msg_to_check_it_0_cnu_68_in_3, msg_to_check_it_0_cnu_68_in_4, msg_to_check_it_0_cnu_68_in_5, msg_to_bit_it_1_vnu_8_in_2, msg_to_bit_it_1_vnu_43_in_2, msg_to_bit_it_1_vnu_82_in_2, msg_to_bit_it_1_vnu_120_in_2, msg_to_bit_it_1_vnu_161_in_2, msg_to_bit_it_1_vnu_197_in_2);
cnu check_node_69_0(msg_to_check_it_0_cnu_69_in_0, msg_to_check_it_0_cnu_69_in_1, msg_to_check_it_0_cnu_69_in_2, msg_to_check_it_0_cnu_69_in_3, msg_to_check_it_0_cnu_69_in_4, msg_to_check_it_0_cnu_69_in_5, msg_to_bit_it_1_vnu_9_in_2, msg_to_bit_it_1_vnu_44_in_2, msg_to_bit_it_1_vnu_83_in_2, msg_to_bit_it_1_vnu_121_in_2, msg_to_bit_it_1_vnu_162_in_2, msg_to_bit_it_1_vnu_165_in_2);
cnu check_node_70_0(msg_to_check_it_0_cnu_70_in_0, msg_to_check_it_0_cnu_70_in_1, msg_to_check_it_0_cnu_70_in_2, msg_to_check_it_0_cnu_70_in_3, msg_to_check_it_0_cnu_70_in_4, msg_to_check_it_0_cnu_70_in_5, msg_to_bit_it_1_vnu_10_in_2, msg_to_bit_it_1_vnu_45_in_2, msg_to_bit_it_1_vnu_84_in_2, msg_to_bit_it_1_vnu_122_in_2, msg_to_bit_it_1_vnu_163_in_2, msg_to_bit_it_1_vnu_166_in_2);
cnu check_node_71_0(msg_to_check_it_0_cnu_71_in_0, msg_to_check_it_0_cnu_71_in_1, msg_to_check_it_0_cnu_71_in_2, msg_to_check_it_0_cnu_71_in_3, msg_to_check_it_0_cnu_71_in_4, msg_to_check_it_0_cnu_71_in_5, msg_to_bit_it_1_vnu_11_in_2, msg_to_bit_it_1_vnu_46_in_2, msg_to_bit_it_1_vnu_85_in_2, msg_to_bit_it_1_vnu_123_in_2, msg_to_bit_it_1_vnu_164_in_2, msg_to_bit_it_1_vnu_167_in_2);
cnu check_node_72_0(msg_to_check_it_0_cnu_72_in_0, msg_to_check_it_0_cnu_72_in_1, msg_to_check_it_0_cnu_72_in_2, msg_to_check_it_0_cnu_72_in_3, msg_to_check_it_0_cnu_72_in_4, msg_to_check_it_0_cnu_72_in_5, msg_to_bit_it_1_vnu_12_in_2, msg_to_bit_it_1_vnu_47_in_2, msg_to_bit_it_1_vnu_86_in_2, msg_to_bit_it_1_vnu_124_in_2, msg_to_bit_it_1_vnu_132_in_2, msg_to_bit_it_1_vnu_168_in_2);
cnu check_node_73_0(msg_to_check_it_0_cnu_73_in_0, msg_to_check_it_0_cnu_73_in_1, msg_to_check_it_0_cnu_73_in_2, msg_to_check_it_0_cnu_73_in_3, msg_to_check_it_0_cnu_73_in_4, msg_to_check_it_0_cnu_73_in_5, msg_to_bit_it_1_vnu_13_in_2, msg_to_bit_it_1_vnu_48_in_2, msg_to_bit_it_1_vnu_87_in_2, msg_to_bit_it_1_vnu_125_in_2, msg_to_bit_it_1_vnu_133_in_2, msg_to_bit_it_1_vnu_169_in_2);
cnu check_node_74_0(msg_to_check_it_0_cnu_74_in_0, msg_to_check_it_0_cnu_74_in_1, msg_to_check_it_0_cnu_74_in_2, msg_to_check_it_0_cnu_74_in_3, msg_to_check_it_0_cnu_74_in_4, msg_to_check_it_0_cnu_74_in_5, msg_to_bit_it_1_vnu_14_in_2, msg_to_bit_it_1_vnu_49_in_2, msg_to_bit_it_1_vnu_88_in_2, msg_to_bit_it_1_vnu_126_in_2, msg_to_bit_it_1_vnu_134_in_2, msg_to_bit_it_1_vnu_170_in_2);
cnu check_node_75_0(msg_to_check_it_0_cnu_75_in_0, msg_to_check_it_0_cnu_75_in_1, msg_to_check_it_0_cnu_75_in_2, msg_to_check_it_0_cnu_75_in_3, msg_to_check_it_0_cnu_75_in_4, msg_to_check_it_0_cnu_75_in_5, msg_to_bit_it_1_vnu_15_in_2, msg_to_bit_it_1_vnu_50_in_2, msg_to_bit_it_1_vnu_89_in_2, msg_to_bit_it_1_vnu_127_in_2, msg_to_bit_it_1_vnu_135_in_2, msg_to_bit_it_1_vnu_171_in_2);
cnu check_node_76_0(msg_to_check_it_0_cnu_76_in_0, msg_to_check_it_0_cnu_76_in_1, msg_to_check_it_0_cnu_76_in_2, msg_to_check_it_0_cnu_76_in_3, msg_to_check_it_0_cnu_76_in_4, msg_to_check_it_0_cnu_76_in_5, msg_to_bit_it_1_vnu_16_in_2, msg_to_bit_it_1_vnu_51_in_2, msg_to_bit_it_1_vnu_90_in_2, msg_to_bit_it_1_vnu_128_in_2, msg_to_bit_it_1_vnu_136_in_2, msg_to_bit_it_1_vnu_172_in_2);
cnu check_node_77_0(msg_to_check_it_0_cnu_77_in_0, msg_to_check_it_0_cnu_77_in_1, msg_to_check_it_0_cnu_77_in_2, msg_to_check_it_0_cnu_77_in_3, msg_to_check_it_0_cnu_77_in_4, msg_to_check_it_0_cnu_77_in_5, msg_to_bit_it_1_vnu_17_in_2, msg_to_bit_it_1_vnu_52_in_2, msg_to_bit_it_1_vnu_91_in_2, msg_to_bit_it_1_vnu_129_in_2, msg_to_bit_it_1_vnu_137_in_2, msg_to_bit_it_1_vnu_173_in_2);
cnu check_node_78_0(msg_to_check_it_0_cnu_78_in_0, msg_to_check_it_0_cnu_78_in_1, msg_to_check_it_0_cnu_78_in_2, msg_to_check_it_0_cnu_78_in_3, msg_to_check_it_0_cnu_78_in_4, msg_to_check_it_0_cnu_78_in_5, msg_to_bit_it_1_vnu_18_in_2, msg_to_bit_it_1_vnu_53_in_2, msg_to_bit_it_1_vnu_92_in_2, msg_to_bit_it_1_vnu_130_in_2, msg_to_bit_it_1_vnu_138_in_2, msg_to_bit_it_1_vnu_174_in_2);
cnu check_node_79_0(msg_to_check_it_0_cnu_79_in_0, msg_to_check_it_0_cnu_79_in_1, msg_to_check_it_0_cnu_79_in_2, msg_to_check_it_0_cnu_79_in_3, msg_to_check_it_0_cnu_79_in_4, msg_to_check_it_0_cnu_79_in_5, msg_to_bit_it_1_vnu_19_in_2, msg_to_bit_it_1_vnu_54_in_2, msg_to_bit_it_1_vnu_93_in_2, msg_to_bit_it_1_vnu_131_in_2, msg_to_bit_it_1_vnu_139_in_2, msg_to_bit_it_1_vnu_175_in_2);
cnu check_node_80_0(msg_to_check_it_0_cnu_80_in_0, msg_to_check_it_0_cnu_80_in_1, msg_to_check_it_0_cnu_80_in_2, msg_to_check_it_0_cnu_80_in_3, msg_to_check_it_0_cnu_80_in_4, msg_to_check_it_0_cnu_80_in_5, msg_to_bit_it_1_vnu_20_in_2, msg_to_bit_it_1_vnu_55_in_2, msg_to_bit_it_1_vnu_94_in_2, msg_to_bit_it_1_vnu_99_in_2, msg_to_bit_it_1_vnu_140_in_2, msg_to_bit_it_1_vnu_176_in_2);
cnu check_node_81_0(msg_to_check_it_0_cnu_81_in_0, msg_to_check_it_0_cnu_81_in_1, msg_to_check_it_0_cnu_81_in_2, msg_to_check_it_0_cnu_81_in_3, msg_to_check_it_0_cnu_81_in_4, msg_to_check_it_0_cnu_81_in_5, msg_to_bit_it_1_vnu_21_in_2, msg_to_bit_it_1_vnu_56_in_2, msg_to_bit_it_1_vnu_95_in_2, msg_to_bit_it_1_vnu_100_in_2, msg_to_bit_it_1_vnu_141_in_2, msg_to_bit_it_1_vnu_177_in_2);
cnu check_node_82_0(msg_to_check_it_0_cnu_82_in_0, msg_to_check_it_0_cnu_82_in_1, msg_to_check_it_0_cnu_82_in_2, msg_to_check_it_0_cnu_82_in_3, msg_to_check_it_0_cnu_82_in_4, msg_to_check_it_0_cnu_82_in_5, msg_to_bit_it_1_vnu_22_in_2, msg_to_bit_it_1_vnu_57_in_2, msg_to_bit_it_1_vnu_96_in_2, msg_to_bit_it_1_vnu_101_in_2, msg_to_bit_it_1_vnu_142_in_2, msg_to_bit_it_1_vnu_178_in_2);
cnu check_node_83_0(msg_to_check_it_0_cnu_83_in_0, msg_to_check_it_0_cnu_83_in_1, msg_to_check_it_0_cnu_83_in_2, msg_to_check_it_0_cnu_83_in_3, msg_to_check_it_0_cnu_83_in_4, msg_to_check_it_0_cnu_83_in_5, msg_to_bit_it_1_vnu_23_in_2, msg_to_bit_it_1_vnu_58_in_2, msg_to_bit_it_1_vnu_97_in_2, msg_to_bit_it_1_vnu_102_in_2, msg_to_bit_it_1_vnu_143_in_2, msg_to_bit_it_1_vnu_179_in_2);
cnu check_node_84_0(msg_to_check_it_0_cnu_84_in_0, msg_to_check_it_0_cnu_84_in_1, msg_to_check_it_0_cnu_84_in_2, msg_to_check_it_0_cnu_84_in_3, msg_to_check_it_0_cnu_84_in_4, msg_to_check_it_0_cnu_84_in_5, msg_to_bit_it_1_vnu_24_in_2, msg_to_bit_it_1_vnu_59_in_2, msg_to_bit_it_1_vnu_98_in_2, msg_to_bit_it_1_vnu_103_in_2, msg_to_bit_it_1_vnu_144_in_2, msg_to_bit_it_1_vnu_180_in_2);
cnu check_node_85_0(msg_to_check_it_0_cnu_85_in_0, msg_to_check_it_0_cnu_85_in_1, msg_to_check_it_0_cnu_85_in_2, msg_to_check_it_0_cnu_85_in_3, msg_to_check_it_0_cnu_85_in_4, msg_to_check_it_0_cnu_85_in_5, msg_to_bit_it_1_vnu_25_in_2, msg_to_bit_it_1_vnu_60_in_2, msg_to_bit_it_1_vnu_66_in_2, msg_to_bit_it_1_vnu_104_in_2, msg_to_bit_it_1_vnu_145_in_2, msg_to_bit_it_1_vnu_181_in_2);
cnu check_node_86_0(msg_to_check_it_0_cnu_86_in_0, msg_to_check_it_0_cnu_86_in_1, msg_to_check_it_0_cnu_86_in_2, msg_to_check_it_0_cnu_86_in_3, msg_to_check_it_0_cnu_86_in_4, msg_to_check_it_0_cnu_86_in_5, msg_to_bit_it_1_vnu_26_in_2, msg_to_bit_it_1_vnu_61_in_2, msg_to_bit_it_1_vnu_67_in_2, msg_to_bit_it_1_vnu_105_in_2, msg_to_bit_it_1_vnu_146_in_2, msg_to_bit_it_1_vnu_182_in_2);
cnu check_node_87_0(msg_to_check_it_0_cnu_87_in_0, msg_to_check_it_0_cnu_87_in_1, msg_to_check_it_0_cnu_87_in_2, msg_to_check_it_0_cnu_87_in_3, msg_to_check_it_0_cnu_87_in_4, msg_to_check_it_0_cnu_87_in_5, msg_to_bit_it_1_vnu_27_in_2, msg_to_bit_it_1_vnu_62_in_2, msg_to_bit_it_1_vnu_68_in_2, msg_to_bit_it_1_vnu_106_in_2, msg_to_bit_it_1_vnu_147_in_2, msg_to_bit_it_1_vnu_183_in_2);
cnu check_node_88_0(msg_to_check_it_0_cnu_88_in_0, msg_to_check_it_0_cnu_88_in_1, msg_to_check_it_0_cnu_88_in_2, msg_to_check_it_0_cnu_88_in_3, msg_to_check_it_0_cnu_88_in_4, msg_to_check_it_0_cnu_88_in_5, msg_to_bit_it_1_vnu_28_in_2, msg_to_bit_it_1_vnu_63_in_2, msg_to_bit_it_1_vnu_69_in_2, msg_to_bit_it_1_vnu_107_in_2, msg_to_bit_it_1_vnu_148_in_2, msg_to_bit_it_1_vnu_184_in_2);
cnu check_node_89_0(msg_to_check_it_0_cnu_89_in_0, msg_to_check_it_0_cnu_89_in_1, msg_to_check_it_0_cnu_89_in_2, msg_to_check_it_0_cnu_89_in_3, msg_to_check_it_0_cnu_89_in_4, msg_to_check_it_0_cnu_89_in_5, msg_to_bit_it_1_vnu_29_in_2, msg_to_bit_it_1_vnu_64_in_2, msg_to_bit_it_1_vnu_70_in_2, msg_to_bit_it_1_vnu_108_in_2, msg_to_bit_it_1_vnu_149_in_2, msg_to_bit_it_1_vnu_185_in_2);
cnu check_node_90_0(msg_to_check_it_0_cnu_90_in_0, msg_to_check_it_0_cnu_90_in_1, msg_to_check_it_0_cnu_90_in_2, msg_to_check_it_0_cnu_90_in_3, msg_to_check_it_0_cnu_90_in_4, msg_to_check_it_0_cnu_90_in_5, msg_to_bit_it_1_vnu_30_in_2, msg_to_bit_it_1_vnu_65_in_2, msg_to_bit_it_1_vnu_71_in_2, msg_to_bit_it_1_vnu_109_in_2, msg_to_bit_it_1_vnu_150_in_2, msg_to_bit_it_1_vnu_186_in_2);
cnu check_node_91_0(msg_to_check_it_0_cnu_91_in_0, msg_to_check_it_0_cnu_91_in_1, msg_to_check_it_0_cnu_91_in_2, msg_to_check_it_0_cnu_91_in_3, msg_to_check_it_0_cnu_91_in_4, msg_to_check_it_0_cnu_91_in_5, msg_to_bit_it_1_vnu_31_in_2, msg_to_bit_it_1_vnu_33_in_2, msg_to_bit_it_1_vnu_72_in_2, msg_to_bit_it_1_vnu_110_in_2, msg_to_bit_it_1_vnu_151_in_2, msg_to_bit_it_1_vnu_187_in_2);
cnu check_node_92_0(msg_to_check_it_0_cnu_92_in_0, msg_to_check_it_0_cnu_92_in_1, msg_to_check_it_0_cnu_92_in_2, msg_to_check_it_0_cnu_92_in_3, msg_to_check_it_0_cnu_92_in_4, msg_to_check_it_0_cnu_92_in_5, msg_to_bit_it_1_vnu_32_in_2, msg_to_bit_it_1_vnu_34_in_2, msg_to_bit_it_1_vnu_73_in_2, msg_to_bit_it_1_vnu_111_in_2, msg_to_bit_it_1_vnu_152_in_2, msg_to_bit_it_1_vnu_188_in_2);
cnu check_node_93_0(msg_to_check_it_0_cnu_93_in_0, msg_to_check_it_0_cnu_93_in_1, msg_to_check_it_0_cnu_93_in_2, msg_to_check_it_0_cnu_93_in_3, msg_to_check_it_0_cnu_93_in_4, msg_to_check_it_0_cnu_93_in_5, msg_to_bit_it_1_vnu_0_in_2, msg_to_bit_it_1_vnu_35_in_2, msg_to_bit_it_1_vnu_74_in_2, msg_to_bit_it_1_vnu_112_in_2, msg_to_bit_it_1_vnu_153_in_2, msg_to_bit_it_1_vnu_189_in_2);
cnu check_node_94_0(msg_to_check_it_0_cnu_94_in_0, msg_to_check_it_0_cnu_94_in_1, msg_to_check_it_0_cnu_94_in_2, msg_to_check_it_0_cnu_94_in_3, msg_to_check_it_0_cnu_94_in_4, msg_to_check_it_0_cnu_94_in_5, msg_to_bit_it_1_vnu_1_in_2, msg_to_bit_it_1_vnu_36_in_2, msg_to_bit_it_1_vnu_75_in_2, msg_to_bit_it_1_vnu_113_in_2, msg_to_bit_it_1_vnu_154_in_2, msg_to_bit_it_1_vnu_190_in_2);
cnu check_node_95_0(msg_to_check_it_0_cnu_95_in_0, msg_to_check_it_0_cnu_95_in_1, msg_to_check_it_0_cnu_95_in_2, msg_to_check_it_0_cnu_95_in_3, msg_to_check_it_0_cnu_95_in_4, msg_to_check_it_0_cnu_95_in_5, msg_to_bit_it_1_vnu_2_in_2, msg_to_bit_it_1_vnu_37_in_2, msg_to_bit_it_1_vnu_76_in_2, msg_to_bit_it_1_vnu_114_in_2, msg_to_bit_it_1_vnu_155_in_2, msg_to_bit_it_1_vnu_191_in_2);
cnu check_node_96_0(msg_to_check_it_0_cnu_96_in_0, msg_to_check_it_0_cnu_96_in_1, msg_to_check_it_0_cnu_96_in_2, msg_to_check_it_0_cnu_96_in_3, msg_to_check_it_0_cnu_96_in_4, msg_to_check_it_0_cnu_96_in_5, msg_to_bit_it_1_vnu_3_in_2, msg_to_bit_it_1_vnu_38_in_2, msg_to_bit_it_1_vnu_77_in_2, msg_to_bit_it_1_vnu_115_in_2, msg_to_bit_it_1_vnu_156_in_2, msg_to_bit_it_1_vnu_192_in_2);
cnu check_node_97_0(msg_to_check_it_0_cnu_97_in_0, msg_to_check_it_0_cnu_97_in_1, msg_to_check_it_0_cnu_97_in_2, msg_to_check_it_0_cnu_97_in_3, msg_to_check_it_0_cnu_97_in_4, msg_to_check_it_0_cnu_97_in_5, msg_to_bit_it_1_vnu_4_in_2, msg_to_bit_it_1_vnu_39_in_2, msg_to_bit_it_1_vnu_78_in_2, msg_to_bit_it_1_vnu_116_in_2, msg_to_bit_it_1_vnu_157_in_2, msg_to_bit_it_1_vnu_193_in_2);
cnu check_node_98_0(msg_to_check_it_0_cnu_98_in_0, msg_to_check_it_0_cnu_98_in_1, msg_to_check_it_0_cnu_98_in_2, msg_to_check_it_0_cnu_98_in_3, msg_to_check_it_0_cnu_98_in_4, msg_to_check_it_0_cnu_98_in_5, msg_to_bit_it_1_vnu_5_in_2, msg_to_bit_it_1_vnu_40_in_2, msg_to_bit_it_1_vnu_79_in_2, msg_to_bit_it_1_vnu_117_in_2, msg_to_bit_it_1_vnu_158_in_2, msg_to_bit_it_1_vnu_194_in_2);


vnu variable_node_0_1(data_0, msg_to_bit_it_1_vnu_0_in_0, msg_to_bit_it_1_vnu_0_in_1, msg_to_bit_it_1_vnu_0_in_2, msg_to_check_it_1_cnu_31_in_0, msg_to_check_it_1_cnu_62_in_0, msg_to_check_it_1_cnu_93_in_0);
vnu variable_node_1_1(data_1, msg_to_bit_it_1_vnu_1_in_0, msg_to_bit_it_1_vnu_1_in_1, msg_to_bit_it_1_vnu_1_in_2, msg_to_check_it_1_cnu_32_in_0, msg_to_check_it_1_cnu_63_in_0, msg_to_check_it_1_cnu_94_in_0);
vnu variable_node_2_1(data_2, msg_to_bit_it_1_vnu_2_in_0, msg_to_bit_it_1_vnu_2_in_1, msg_to_bit_it_1_vnu_2_in_2, msg_to_check_it_1_cnu_0_in_0, msg_to_check_it_1_cnu_64_in_0, msg_to_check_it_1_cnu_95_in_0);
vnu variable_node_3_1(data_3, msg_to_bit_it_1_vnu_3_in_0, msg_to_bit_it_1_vnu_3_in_1, msg_to_bit_it_1_vnu_3_in_2, msg_to_check_it_1_cnu_1_in_0, msg_to_check_it_1_cnu_65_in_0, msg_to_check_it_1_cnu_96_in_0);
vnu variable_node_4_1(data_4, msg_to_bit_it_1_vnu_4_in_0, msg_to_bit_it_1_vnu_4_in_1, msg_to_bit_it_1_vnu_4_in_2, msg_to_check_it_1_cnu_2_in_0, msg_to_check_it_1_cnu_33_in_0, msg_to_check_it_1_cnu_97_in_0);
vnu variable_node_5_1(data_5, msg_to_bit_it_1_vnu_5_in_0, msg_to_bit_it_1_vnu_5_in_1, msg_to_bit_it_1_vnu_5_in_2, msg_to_check_it_1_cnu_3_in_0, msg_to_check_it_1_cnu_34_in_0, msg_to_check_it_1_cnu_98_in_0);
vnu variable_node_6_1(data_6, msg_to_bit_it_1_vnu_6_in_0, msg_to_bit_it_1_vnu_6_in_1, msg_to_bit_it_1_vnu_6_in_2, msg_to_check_it_1_cnu_4_in_0, msg_to_check_it_1_cnu_35_in_0, msg_to_check_it_1_cnu_66_in_0);
vnu variable_node_7_1(data_7, msg_to_bit_it_1_vnu_7_in_0, msg_to_bit_it_1_vnu_7_in_1, msg_to_bit_it_1_vnu_7_in_2, msg_to_check_it_1_cnu_5_in_0, msg_to_check_it_1_cnu_36_in_0, msg_to_check_it_1_cnu_67_in_0);
vnu variable_node_8_1(data_8, msg_to_bit_it_1_vnu_8_in_0, msg_to_bit_it_1_vnu_8_in_1, msg_to_bit_it_1_vnu_8_in_2, msg_to_check_it_1_cnu_6_in_0, msg_to_check_it_1_cnu_37_in_0, msg_to_check_it_1_cnu_68_in_0);
vnu variable_node_9_1(data_9, msg_to_bit_it_1_vnu_9_in_0, msg_to_bit_it_1_vnu_9_in_1, msg_to_bit_it_1_vnu_9_in_2, msg_to_check_it_1_cnu_7_in_0, msg_to_check_it_1_cnu_38_in_0, msg_to_check_it_1_cnu_69_in_0);
vnu variable_node_10_1(data_10, msg_to_bit_it_1_vnu_10_in_0, msg_to_bit_it_1_vnu_10_in_1, msg_to_bit_it_1_vnu_10_in_2, msg_to_check_it_1_cnu_8_in_0, msg_to_check_it_1_cnu_39_in_0, msg_to_check_it_1_cnu_70_in_0);
vnu variable_node_11_1(data_11, msg_to_bit_it_1_vnu_11_in_0, msg_to_bit_it_1_vnu_11_in_1, msg_to_bit_it_1_vnu_11_in_2, msg_to_check_it_1_cnu_9_in_0, msg_to_check_it_1_cnu_40_in_0, msg_to_check_it_1_cnu_71_in_0);
vnu variable_node_12_1(data_12, msg_to_bit_it_1_vnu_12_in_0, msg_to_bit_it_1_vnu_12_in_1, msg_to_bit_it_1_vnu_12_in_2, msg_to_check_it_1_cnu_10_in_0, msg_to_check_it_1_cnu_41_in_0, msg_to_check_it_1_cnu_72_in_0);
vnu variable_node_13_1(data_13, msg_to_bit_it_1_vnu_13_in_0, msg_to_bit_it_1_vnu_13_in_1, msg_to_bit_it_1_vnu_13_in_2, msg_to_check_it_1_cnu_11_in_0, msg_to_check_it_1_cnu_42_in_0, msg_to_check_it_1_cnu_73_in_0);
vnu variable_node_14_1(data_14, msg_to_bit_it_1_vnu_14_in_0, msg_to_bit_it_1_vnu_14_in_1, msg_to_bit_it_1_vnu_14_in_2, msg_to_check_it_1_cnu_12_in_0, msg_to_check_it_1_cnu_43_in_0, msg_to_check_it_1_cnu_74_in_0);
vnu variable_node_15_1(data_15, msg_to_bit_it_1_vnu_15_in_0, msg_to_bit_it_1_vnu_15_in_1, msg_to_bit_it_1_vnu_15_in_2, msg_to_check_it_1_cnu_13_in_0, msg_to_check_it_1_cnu_44_in_0, msg_to_check_it_1_cnu_75_in_0);
vnu variable_node_16_1(data_16, msg_to_bit_it_1_vnu_16_in_0, msg_to_bit_it_1_vnu_16_in_1, msg_to_bit_it_1_vnu_16_in_2, msg_to_check_it_1_cnu_14_in_0, msg_to_check_it_1_cnu_45_in_0, msg_to_check_it_1_cnu_76_in_0);
vnu variable_node_17_1(data_17, msg_to_bit_it_1_vnu_17_in_0, msg_to_bit_it_1_vnu_17_in_1, msg_to_bit_it_1_vnu_17_in_2, msg_to_check_it_1_cnu_15_in_0, msg_to_check_it_1_cnu_46_in_0, msg_to_check_it_1_cnu_77_in_0);
vnu variable_node_18_1(data_18, msg_to_bit_it_1_vnu_18_in_0, msg_to_bit_it_1_vnu_18_in_1, msg_to_bit_it_1_vnu_18_in_2, msg_to_check_it_1_cnu_16_in_0, msg_to_check_it_1_cnu_47_in_0, msg_to_check_it_1_cnu_78_in_0);
vnu variable_node_19_1(data_19, msg_to_bit_it_1_vnu_19_in_0, msg_to_bit_it_1_vnu_19_in_1, msg_to_bit_it_1_vnu_19_in_2, msg_to_check_it_1_cnu_17_in_0, msg_to_check_it_1_cnu_48_in_0, msg_to_check_it_1_cnu_79_in_0);
vnu variable_node_20_1(data_20, msg_to_bit_it_1_vnu_20_in_0, msg_to_bit_it_1_vnu_20_in_1, msg_to_bit_it_1_vnu_20_in_2, msg_to_check_it_1_cnu_18_in_0, msg_to_check_it_1_cnu_49_in_0, msg_to_check_it_1_cnu_80_in_0);
vnu variable_node_21_1(data_21, msg_to_bit_it_1_vnu_21_in_0, msg_to_bit_it_1_vnu_21_in_1, msg_to_bit_it_1_vnu_21_in_2, msg_to_check_it_1_cnu_19_in_0, msg_to_check_it_1_cnu_50_in_0, msg_to_check_it_1_cnu_81_in_0);
vnu variable_node_22_1(data_22, msg_to_bit_it_1_vnu_22_in_0, msg_to_bit_it_1_vnu_22_in_1, msg_to_bit_it_1_vnu_22_in_2, msg_to_check_it_1_cnu_20_in_0, msg_to_check_it_1_cnu_51_in_0, msg_to_check_it_1_cnu_82_in_0);
vnu variable_node_23_1(data_23, msg_to_bit_it_1_vnu_23_in_0, msg_to_bit_it_1_vnu_23_in_1, msg_to_bit_it_1_vnu_23_in_2, msg_to_check_it_1_cnu_21_in_0, msg_to_check_it_1_cnu_52_in_0, msg_to_check_it_1_cnu_83_in_0);
vnu variable_node_24_1(data_24, msg_to_bit_it_1_vnu_24_in_0, msg_to_bit_it_1_vnu_24_in_1, msg_to_bit_it_1_vnu_24_in_2, msg_to_check_it_1_cnu_22_in_0, msg_to_check_it_1_cnu_53_in_0, msg_to_check_it_1_cnu_84_in_0);
vnu variable_node_25_1(data_25, msg_to_bit_it_1_vnu_25_in_0, msg_to_bit_it_1_vnu_25_in_1, msg_to_bit_it_1_vnu_25_in_2, msg_to_check_it_1_cnu_23_in_0, msg_to_check_it_1_cnu_54_in_0, msg_to_check_it_1_cnu_85_in_0);
vnu variable_node_26_1(data_26, msg_to_bit_it_1_vnu_26_in_0, msg_to_bit_it_1_vnu_26_in_1, msg_to_bit_it_1_vnu_26_in_2, msg_to_check_it_1_cnu_24_in_0, msg_to_check_it_1_cnu_55_in_0, msg_to_check_it_1_cnu_86_in_0);
vnu variable_node_27_1(data_27, msg_to_bit_it_1_vnu_27_in_0, msg_to_bit_it_1_vnu_27_in_1, msg_to_bit_it_1_vnu_27_in_2, msg_to_check_it_1_cnu_25_in_0, msg_to_check_it_1_cnu_56_in_0, msg_to_check_it_1_cnu_87_in_0);
vnu variable_node_28_1(data_28, msg_to_bit_it_1_vnu_28_in_0, msg_to_bit_it_1_vnu_28_in_1, msg_to_bit_it_1_vnu_28_in_2, msg_to_check_it_1_cnu_26_in_0, msg_to_check_it_1_cnu_57_in_0, msg_to_check_it_1_cnu_88_in_0);
vnu variable_node_29_1(data_29, msg_to_bit_it_1_vnu_29_in_0, msg_to_bit_it_1_vnu_29_in_1, msg_to_bit_it_1_vnu_29_in_2, msg_to_check_it_1_cnu_27_in_0, msg_to_check_it_1_cnu_58_in_0, msg_to_check_it_1_cnu_89_in_0);
vnu variable_node_30_1(data_30, msg_to_bit_it_1_vnu_30_in_0, msg_to_bit_it_1_vnu_30_in_1, msg_to_bit_it_1_vnu_30_in_2, msg_to_check_it_1_cnu_28_in_0, msg_to_check_it_1_cnu_59_in_0, msg_to_check_it_1_cnu_90_in_0);
vnu variable_node_31_1(data_31, msg_to_bit_it_1_vnu_31_in_0, msg_to_bit_it_1_vnu_31_in_1, msg_to_bit_it_1_vnu_31_in_2, msg_to_check_it_1_cnu_29_in_0, msg_to_check_it_1_cnu_60_in_0, msg_to_check_it_1_cnu_91_in_0);
vnu variable_node_32_1(data_32, msg_to_bit_it_1_vnu_32_in_0, msg_to_bit_it_1_vnu_32_in_1, msg_to_bit_it_1_vnu_32_in_2, msg_to_check_it_1_cnu_30_in_0, msg_to_check_it_1_cnu_61_in_0, msg_to_check_it_1_cnu_92_in_0);
vnu variable_node_33_1(data_33, msg_to_bit_it_1_vnu_33_in_0, msg_to_bit_it_1_vnu_33_in_1, msg_to_bit_it_1_vnu_33_in_2, msg_to_check_it_1_cnu_30_in_1, msg_to_check_it_1_cnu_61_in_1, msg_to_check_it_1_cnu_91_in_1);
vnu variable_node_34_1(data_34, msg_to_bit_it_1_vnu_34_in_0, msg_to_bit_it_1_vnu_34_in_1, msg_to_bit_it_1_vnu_34_in_2, msg_to_check_it_1_cnu_31_in_1, msg_to_check_it_1_cnu_62_in_1, msg_to_check_it_1_cnu_92_in_1);
vnu variable_node_35_1(data_35, msg_to_bit_it_1_vnu_35_in_0, msg_to_bit_it_1_vnu_35_in_1, msg_to_bit_it_1_vnu_35_in_2, msg_to_check_it_1_cnu_32_in_1, msg_to_check_it_1_cnu_63_in_1, msg_to_check_it_1_cnu_93_in_1);
vnu variable_node_36_1(data_36, msg_to_bit_it_1_vnu_36_in_0, msg_to_bit_it_1_vnu_36_in_1, msg_to_bit_it_1_vnu_36_in_2, msg_to_check_it_1_cnu_0_in_1, msg_to_check_it_1_cnu_64_in_1, msg_to_check_it_1_cnu_94_in_1);
vnu variable_node_37_1(data_37, msg_to_bit_it_1_vnu_37_in_0, msg_to_bit_it_1_vnu_37_in_1, msg_to_bit_it_1_vnu_37_in_2, msg_to_check_it_1_cnu_1_in_1, msg_to_check_it_1_cnu_65_in_1, msg_to_check_it_1_cnu_95_in_1);
vnu variable_node_38_1(data_38, msg_to_bit_it_1_vnu_38_in_0, msg_to_bit_it_1_vnu_38_in_1, msg_to_bit_it_1_vnu_38_in_2, msg_to_check_it_1_cnu_2_in_1, msg_to_check_it_1_cnu_33_in_1, msg_to_check_it_1_cnu_96_in_1);
vnu variable_node_39_1(data_39, msg_to_bit_it_1_vnu_39_in_0, msg_to_bit_it_1_vnu_39_in_1, msg_to_bit_it_1_vnu_39_in_2, msg_to_check_it_1_cnu_3_in_1, msg_to_check_it_1_cnu_34_in_1, msg_to_check_it_1_cnu_97_in_1);
vnu variable_node_40_1(data_40, msg_to_bit_it_1_vnu_40_in_0, msg_to_bit_it_1_vnu_40_in_1, msg_to_bit_it_1_vnu_40_in_2, msg_to_check_it_1_cnu_4_in_1, msg_to_check_it_1_cnu_35_in_1, msg_to_check_it_1_cnu_98_in_1);
vnu variable_node_41_1(data_41, msg_to_bit_it_1_vnu_41_in_0, msg_to_bit_it_1_vnu_41_in_1, msg_to_bit_it_1_vnu_41_in_2, msg_to_check_it_1_cnu_5_in_1, msg_to_check_it_1_cnu_36_in_1, msg_to_check_it_1_cnu_66_in_1);
vnu variable_node_42_1(data_42, msg_to_bit_it_1_vnu_42_in_0, msg_to_bit_it_1_vnu_42_in_1, msg_to_bit_it_1_vnu_42_in_2, msg_to_check_it_1_cnu_6_in_1, msg_to_check_it_1_cnu_37_in_1, msg_to_check_it_1_cnu_67_in_1);
vnu variable_node_43_1(data_43, msg_to_bit_it_1_vnu_43_in_0, msg_to_bit_it_1_vnu_43_in_1, msg_to_bit_it_1_vnu_43_in_2, msg_to_check_it_1_cnu_7_in_1, msg_to_check_it_1_cnu_38_in_1, msg_to_check_it_1_cnu_68_in_1);
vnu variable_node_44_1(data_44, msg_to_bit_it_1_vnu_44_in_0, msg_to_bit_it_1_vnu_44_in_1, msg_to_bit_it_1_vnu_44_in_2, msg_to_check_it_1_cnu_8_in_1, msg_to_check_it_1_cnu_39_in_1, msg_to_check_it_1_cnu_69_in_1);
vnu variable_node_45_1(data_45, msg_to_bit_it_1_vnu_45_in_0, msg_to_bit_it_1_vnu_45_in_1, msg_to_bit_it_1_vnu_45_in_2, msg_to_check_it_1_cnu_9_in_1, msg_to_check_it_1_cnu_40_in_1, msg_to_check_it_1_cnu_70_in_1);
vnu variable_node_46_1(data_46, msg_to_bit_it_1_vnu_46_in_0, msg_to_bit_it_1_vnu_46_in_1, msg_to_bit_it_1_vnu_46_in_2, msg_to_check_it_1_cnu_10_in_1, msg_to_check_it_1_cnu_41_in_1, msg_to_check_it_1_cnu_71_in_1);
vnu variable_node_47_1(data_47, msg_to_bit_it_1_vnu_47_in_0, msg_to_bit_it_1_vnu_47_in_1, msg_to_bit_it_1_vnu_47_in_2, msg_to_check_it_1_cnu_11_in_1, msg_to_check_it_1_cnu_42_in_1, msg_to_check_it_1_cnu_72_in_1);
vnu variable_node_48_1(data_48, msg_to_bit_it_1_vnu_48_in_0, msg_to_bit_it_1_vnu_48_in_1, msg_to_bit_it_1_vnu_48_in_2, msg_to_check_it_1_cnu_12_in_1, msg_to_check_it_1_cnu_43_in_1, msg_to_check_it_1_cnu_73_in_1);
vnu variable_node_49_1(data_49, msg_to_bit_it_1_vnu_49_in_0, msg_to_bit_it_1_vnu_49_in_1, msg_to_bit_it_1_vnu_49_in_2, msg_to_check_it_1_cnu_13_in_1, msg_to_check_it_1_cnu_44_in_1, msg_to_check_it_1_cnu_74_in_1);
vnu variable_node_50_1(data_50, msg_to_bit_it_1_vnu_50_in_0, msg_to_bit_it_1_vnu_50_in_1, msg_to_bit_it_1_vnu_50_in_2, msg_to_check_it_1_cnu_14_in_1, msg_to_check_it_1_cnu_45_in_1, msg_to_check_it_1_cnu_75_in_1);
vnu variable_node_51_1(data_51, msg_to_bit_it_1_vnu_51_in_0, msg_to_bit_it_1_vnu_51_in_1, msg_to_bit_it_1_vnu_51_in_2, msg_to_check_it_1_cnu_15_in_1, msg_to_check_it_1_cnu_46_in_1, msg_to_check_it_1_cnu_76_in_1);
vnu variable_node_52_1(data_52, msg_to_bit_it_1_vnu_52_in_0, msg_to_bit_it_1_vnu_52_in_1, msg_to_bit_it_1_vnu_52_in_2, msg_to_check_it_1_cnu_16_in_1, msg_to_check_it_1_cnu_47_in_1, msg_to_check_it_1_cnu_77_in_1);
vnu variable_node_53_1(data_53, msg_to_bit_it_1_vnu_53_in_0, msg_to_bit_it_1_vnu_53_in_1, msg_to_bit_it_1_vnu_53_in_2, msg_to_check_it_1_cnu_17_in_1, msg_to_check_it_1_cnu_48_in_1, msg_to_check_it_1_cnu_78_in_1);
vnu variable_node_54_1(data_54, msg_to_bit_it_1_vnu_54_in_0, msg_to_bit_it_1_vnu_54_in_1, msg_to_bit_it_1_vnu_54_in_2, msg_to_check_it_1_cnu_18_in_1, msg_to_check_it_1_cnu_49_in_1, msg_to_check_it_1_cnu_79_in_1);
vnu variable_node_55_1(data_55, msg_to_bit_it_1_vnu_55_in_0, msg_to_bit_it_1_vnu_55_in_1, msg_to_bit_it_1_vnu_55_in_2, msg_to_check_it_1_cnu_19_in_1, msg_to_check_it_1_cnu_50_in_1, msg_to_check_it_1_cnu_80_in_1);
vnu variable_node_56_1(data_56, msg_to_bit_it_1_vnu_56_in_0, msg_to_bit_it_1_vnu_56_in_1, msg_to_bit_it_1_vnu_56_in_2, msg_to_check_it_1_cnu_20_in_1, msg_to_check_it_1_cnu_51_in_1, msg_to_check_it_1_cnu_81_in_1);
vnu variable_node_57_1(data_57, msg_to_bit_it_1_vnu_57_in_0, msg_to_bit_it_1_vnu_57_in_1, msg_to_bit_it_1_vnu_57_in_2, msg_to_check_it_1_cnu_21_in_1, msg_to_check_it_1_cnu_52_in_1, msg_to_check_it_1_cnu_82_in_1);
vnu variable_node_58_1(data_58, msg_to_bit_it_1_vnu_58_in_0, msg_to_bit_it_1_vnu_58_in_1, msg_to_bit_it_1_vnu_58_in_2, msg_to_check_it_1_cnu_22_in_1, msg_to_check_it_1_cnu_53_in_1, msg_to_check_it_1_cnu_83_in_1);
vnu variable_node_59_1(data_59, msg_to_bit_it_1_vnu_59_in_0, msg_to_bit_it_1_vnu_59_in_1, msg_to_bit_it_1_vnu_59_in_2, msg_to_check_it_1_cnu_23_in_1, msg_to_check_it_1_cnu_54_in_1, msg_to_check_it_1_cnu_84_in_1);
vnu variable_node_60_1(data_60, msg_to_bit_it_1_vnu_60_in_0, msg_to_bit_it_1_vnu_60_in_1, msg_to_bit_it_1_vnu_60_in_2, msg_to_check_it_1_cnu_24_in_1, msg_to_check_it_1_cnu_55_in_1, msg_to_check_it_1_cnu_85_in_1);
vnu variable_node_61_1(data_61, msg_to_bit_it_1_vnu_61_in_0, msg_to_bit_it_1_vnu_61_in_1, msg_to_bit_it_1_vnu_61_in_2, msg_to_check_it_1_cnu_25_in_1, msg_to_check_it_1_cnu_56_in_1, msg_to_check_it_1_cnu_86_in_1);
vnu variable_node_62_1(data_62, msg_to_bit_it_1_vnu_62_in_0, msg_to_bit_it_1_vnu_62_in_1, msg_to_bit_it_1_vnu_62_in_2, msg_to_check_it_1_cnu_26_in_1, msg_to_check_it_1_cnu_57_in_1, msg_to_check_it_1_cnu_87_in_1);
vnu variable_node_63_1(data_63, msg_to_bit_it_1_vnu_63_in_0, msg_to_bit_it_1_vnu_63_in_1, msg_to_bit_it_1_vnu_63_in_2, msg_to_check_it_1_cnu_27_in_1, msg_to_check_it_1_cnu_58_in_1, msg_to_check_it_1_cnu_88_in_1);
vnu variable_node_64_1(data_64, msg_to_bit_it_1_vnu_64_in_0, msg_to_bit_it_1_vnu_64_in_1, msg_to_bit_it_1_vnu_64_in_2, msg_to_check_it_1_cnu_28_in_1, msg_to_check_it_1_cnu_59_in_1, msg_to_check_it_1_cnu_89_in_1);
vnu variable_node_65_1(data_65, msg_to_bit_it_1_vnu_65_in_0, msg_to_bit_it_1_vnu_65_in_1, msg_to_bit_it_1_vnu_65_in_2, msg_to_check_it_1_cnu_29_in_1, msg_to_check_it_1_cnu_60_in_1, msg_to_check_it_1_cnu_90_in_1);
vnu variable_node_66_1(data_66, msg_to_bit_it_1_vnu_66_in_0, msg_to_bit_it_1_vnu_66_in_1, msg_to_bit_it_1_vnu_66_in_2, msg_to_check_it_1_cnu_26_in_2, msg_to_check_it_1_cnu_55_in_2, msg_to_check_it_1_cnu_85_in_2);
vnu variable_node_67_1(data_67, msg_to_bit_it_1_vnu_67_in_0, msg_to_bit_it_1_vnu_67_in_1, msg_to_bit_it_1_vnu_67_in_2, msg_to_check_it_1_cnu_27_in_2, msg_to_check_it_1_cnu_56_in_2, msg_to_check_it_1_cnu_86_in_2);
vnu variable_node_68_1(data_68, msg_to_bit_it_1_vnu_68_in_0, msg_to_bit_it_1_vnu_68_in_1, msg_to_bit_it_1_vnu_68_in_2, msg_to_check_it_1_cnu_28_in_2, msg_to_check_it_1_cnu_57_in_2, msg_to_check_it_1_cnu_87_in_2);
vnu variable_node_69_1(data_69, msg_to_bit_it_1_vnu_69_in_0, msg_to_bit_it_1_vnu_69_in_1, msg_to_bit_it_1_vnu_69_in_2, msg_to_check_it_1_cnu_29_in_2, msg_to_check_it_1_cnu_58_in_2, msg_to_check_it_1_cnu_88_in_2);
vnu variable_node_70_1(data_70, msg_to_bit_it_1_vnu_70_in_0, msg_to_bit_it_1_vnu_70_in_1, msg_to_bit_it_1_vnu_70_in_2, msg_to_check_it_1_cnu_30_in_2, msg_to_check_it_1_cnu_59_in_2, msg_to_check_it_1_cnu_89_in_2);
vnu variable_node_71_1(data_71, msg_to_bit_it_1_vnu_71_in_0, msg_to_bit_it_1_vnu_71_in_1, msg_to_bit_it_1_vnu_71_in_2, msg_to_check_it_1_cnu_31_in_2, msg_to_check_it_1_cnu_60_in_2, msg_to_check_it_1_cnu_90_in_2);
vnu variable_node_72_1(data_72, msg_to_bit_it_1_vnu_72_in_0, msg_to_bit_it_1_vnu_72_in_1, msg_to_bit_it_1_vnu_72_in_2, msg_to_check_it_1_cnu_32_in_2, msg_to_check_it_1_cnu_61_in_2, msg_to_check_it_1_cnu_91_in_2);
vnu variable_node_73_1(data_73, msg_to_bit_it_1_vnu_73_in_0, msg_to_bit_it_1_vnu_73_in_1, msg_to_bit_it_1_vnu_73_in_2, msg_to_check_it_1_cnu_0_in_2, msg_to_check_it_1_cnu_62_in_2, msg_to_check_it_1_cnu_92_in_2);
vnu variable_node_74_1(data_74, msg_to_bit_it_1_vnu_74_in_0, msg_to_bit_it_1_vnu_74_in_1, msg_to_bit_it_1_vnu_74_in_2, msg_to_check_it_1_cnu_1_in_2, msg_to_check_it_1_cnu_63_in_2, msg_to_check_it_1_cnu_93_in_2);
vnu variable_node_75_1(data_75, msg_to_bit_it_1_vnu_75_in_0, msg_to_bit_it_1_vnu_75_in_1, msg_to_bit_it_1_vnu_75_in_2, msg_to_check_it_1_cnu_2_in_2, msg_to_check_it_1_cnu_64_in_2, msg_to_check_it_1_cnu_94_in_2);
vnu variable_node_76_1(data_76, msg_to_bit_it_1_vnu_76_in_0, msg_to_bit_it_1_vnu_76_in_1, msg_to_bit_it_1_vnu_76_in_2, msg_to_check_it_1_cnu_3_in_2, msg_to_check_it_1_cnu_65_in_2, msg_to_check_it_1_cnu_95_in_2);
vnu variable_node_77_1(data_77, msg_to_bit_it_1_vnu_77_in_0, msg_to_bit_it_1_vnu_77_in_1, msg_to_bit_it_1_vnu_77_in_2, msg_to_check_it_1_cnu_4_in_2, msg_to_check_it_1_cnu_33_in_2, msg_to_check_it_1_cnu_96_in_2);
vnu variable_node_78_1(data_78, msg_to_bit_it_1_vnu_78_in_0, msg_to_bit_it_1_vnu_78_in_1, msg_to_bit_it_1_vnu_78_in_2, msg_to_check_it_1_cnu_5_in_2, msg_to_check_it_1_cnu_34_in_2, msg_to_check_it_1_cnu_97_in_2);
vnu variable_node_79_1(data_79, msg_to_bit_it_1_vnu_79_in_0, msg_to_bit_it_1_vnu_79_in_1, msg_to_bit_it_1_vnu_79_in_2, msg_to_check_it_1_cnu_6_in_2, msg_to_check_it_1_cnu_35_in_2, msg_to_check_it_1_cnu_98_in_2);
vnu variable_node_80_1(data_80, msg_to_bit_it_1_vnu_80_in_0, msg_to_bit_it_1_vnu_80_in_1, msg_to_bit_it_1_vnu_80_in_2, msg_to_check_it_1_cnu_7_in_2, msg_to_check_it_1_cnu_36_in_2, msg_to_check_it_1_cnu_66_in_2);
vnu variable_node_81_1(data_81, msg_to_bit_it_1_vnu_81_in_0, msg_to_bit_it_1_vnu_81_in_1, msg_to_bit_it_1_vnu_81_in_2, msg_to_check_it_1_cnu_8_in_2, msg_to_check_it_1_cnu_37_in_2, msg_to_check_it_1_cnu_67_in_2);
vnu variable_node_82_1(data_82, msg_to_bit_it_1_vnu_82_in_0, msg_to_bit_it_1_vnu_82_in_1, msg_to_bit_it_1_vnu_82_in_2, msg_to_check_it_1_cnu_9_in_2, msg_to_check_it_1_cnu_38_in_2, msg_to_check_it_1_cnu_68_in_2);
vnu variable_node_83_1(data_83, msg_to_bit_it_1_vnu_83_in_0, msg_to_bit_it_1_vnu_83_in_1, msg_to_bit_it_1_vnu_83_in_2, msg_to_check_it_1_cnu_10_in_2, msg_to_check_it_1_cnu_39_in_2, msg_to_check_it_1_cnu_69_in_2);
vnu variable_node_84_1(data_84, msg_to_bit_it_1_vnu_84_in_0, msg_to_bit_it_1_vnu_84_in_1, msg_to_bit_it_1_vnu_84_in_2, msg_to_check_it_1_cnu_11_in_2, msg_to_check_it_1_cnu_40_in_2, msg_to_check_it_1_cnu_70_in_2);
vnu variable_node_85_1(data_85, msg_to_bit_it_1_vnu_85_in_0, msg_to_bit_it_1_vnu_85_in_1, msg_to_bit_it_1_vnu_85_in_2, msg_to_check_it_1_cnu_12_in_2, msg_to_check_it_1_cnu_41_in_2, msg_to_check_it_1_cnu_71_in_2);
vnu variable_node_86_1(data_86, msg_to_bit_it_1_vnu_86_in_0, msg_to_bit_it_1_vnu_86_in_1, msg_to_bit_it_1_vnu_86_in_2, msg_to_check_it_1_cnu_13_in_2, msg_to_check_it_1_cnu_42_in_2, msg_to_check_it_1_cnu_72_in_2);
vnu variable_node_87_1(data_87, msg_to_bit_it_1_vnu_87_in_0, msg_to_bit_it_1_vnu_87_in_1, msg_to_bit_it_1_vnu_87_in_2, msg_to_check_it_1_cnu_14_in_2, msg_to_check_it_1_cnu_43_in_2, msg_to_check_it_1_cnu_73_in_2);
vnu variable_node_88_1(data_88, msg_to_bit_it_1_vnu_88_in_0, msg_to_bit_it_1_vnu_88_in_1, msg_to_bit_it_1_vnu_88_in_2, msg_to_check_it_1_cnu_15_in_2, msg_to_check_it_1_cnu_44_in_2, msg_to_check_it_1_cnu_74_in_2);
vnu variable_node_89_1(data_89, msg_to_bit_it_1_vnu_89_in_0, msg_to_bit_it_1_vnu_89_in_1, msg_to_bit_it_1_vnu_89_in_2, msg_to_check_it_1_cnu_16_in_2, msg_to_check_it_1_cnu_45_in_2, msg_to_check_it_1_cnu_75_in_2);
vnu variable_node_90_1(data_90, msg_to_bit_it_1_vnu_90_in_0, msg_to_bit_it_1_vnu_90_in_1, msg_to_bit_it_1_vnu_90_in_2, msg_to_check_it_1_cnu_17_in_2, msg_to_check_it_1_cnu_46_in_2, msg_to_check_it_1_cnu_76_in_2);
vnu variable_node_91_1(data_91, msg_to_bit_it_1_vnu_91_in_0, msg_to_bit_it_1_vnu_91_in_1, msg_to_bit_it_1_vnu_91_in_2, msg_to_check_it_1_cnu_18_in_2, msg_to_check_it_1_cnu_47_in_2, msg_to_check_it_1_cnu_77_in_2);
vnu variable_node_92_1(data_92, msg_to_bit_it_1_vnu_92_in_0, msg_to_bit_it_1_vnu_92_in_1, msg_to_bit_it_1_vnu_92_in_2, msg_to_check_it_1_cnu_19_in_2, msg_to_check_it_1_cnu_48_in_2, msg_to_check_it_1_cnu_78_in_2);
vnu variable_node_93_1(data_93, msg_to_bit_it_1_vnu_93_in_0, msg_to_bit_it_1_vnu_93_in_1, msg_to_bit_it_1_vnu_93_in_2, msg_to_check_it_1_cnu_20_in_2, msg_to_check_it_1_cnu_49_in_2, msg_to_check_it_1_cnu_79_in_2);
vnu variable_node_94_1(data_94, msg_to_bit_it_1_vnu_94_in_0, msg_to_bit_it_1_vnu_94_in_1, msg_to_bit_it_1_vnu_94_in_2, msg_to_check_it_1_cnu_21_in_2, msg_to_check_it_1_cnu_50_in_2, msg_to_check_it_1_cnu_80_in_2);
vnu variable_node_95_1(data_95, msg_to_bit_it_1_vnu_95_in_0, msg_to_bit_it_1_vnu_95_in_1, msg_to_bit_it_1_vnu_95_in_2, msg_to_check_it_1_cnu_22_in_2, msg_to_check_it_1_cnu_51_in_2, msg_to_check_it_1_cnu_81_in_2);
vnu variable_node_96_1(data_96, msg_to_bit_it_1_vnu_96_in_0, msg_to_bit_it_1_vnu_96_in_1, msg_to_bit_it_1_vnu_96_in_2, msg_to_check_it_1_cnu_23_in_2, msg_to_check_it_1_cnu_52_in_2, msg_to_check_it_1_cnu_82_in_2);
vnu variable_node_97_1(data_97, msg_to_bit_it_1_vnu_97_in_0, msg_to_bit_it_1_vnu_97_in_1, msg_to_bit_it_1_vnu_97_in_2, msg_to_check_it_1_cnu_24_in_2, msg_to_check_it_1_cnu_53_in_2, msg_to_check_it_1_cnu_83_in_2);
vnu variable_node_98_1(data_98, msg_to_bit_it_1_vnu_98_in_0, msg_to_bit_it_1_vnu_98_in_1, msg_to_bit_it_1_vnu_98_in_2, msg_to_check_it_1_cnu_25_in_2, msg_to_check_it_1_cnu_54_in_2, msg_to_check_it_1_cnu_84_in_2);
vnu variable_node_99_1(data_99, msg_to_bit_it_1_vnu_99_in_0, msg_to_bit_it_1_vnu_99_in_1, msg_to_bit_it_1_vnu_99_in_2, msg_to_check_it_1_cnu_24_in_3, msg_to_check_it_1_cnu_54_in_3, msg_to_check_it_1_cnu_80_in_3);
vnu variable_node_100_1(data_100, msg_to_bit_it_1_vnu_100_in_0, msg_to_bit_it_1_vnu_100_in_1, msg_to_bit_it_1_vnu_100_in_2, msg_to_check_it_1_cnu_25_in_3, msg_to_check_it_1_cnu_55_in_3, msg_to_check_it_1_cnu_81_in_3);
vnu variable_node_101_1(data_101, msg_to_bit_it_1_vnu_101_in_0, msg_to_bit_it_1_vnu_101_in_1, msg_to_bit_it_1_vnu_101_in_2, msg_to_check_it_1_cnu_26_in_3, msg_to_check_it_1_cnu_56_in_3, msg_to_check_it_1_cnu_82_in_3);
vnu variable_node_102_1(data_102, msg_to_bit_it_1_vnu_102_in_0, msg_to_bit_it_1_vnu_102_in_1, msg_to_bit_it_1_vnu_102_in_2, msg_to_check_it_1_cnu_27_in_3, msg_to_check_it_1_cnu_57_in_3, msg_to_check_it_1_cnu_83_in_3);
vnu variable_node_103_1(data_103, msg_to_bit_it_1_vnu_103_in_0, msg_to_bit_it_1_vnu_103_in_1, msg_to_bit_it_1_vnu_103_in_2, msg_to_check_it_1_cnu_28_in_3, msg_to_check_it_1_cnu_58_in_3, msg_to_check_it_1_cnu_84_in_3);
vnu variable_node_104_1(data_104, msg_to_bit_it_1_vnu_104_in_0, msg_to_bit_it_1_vnu_104_in_1, msg_to_bit_it_1_vnu_104_in_2, msg_to_check_it_1_cnu_29_in_3, msg_to_check_it_1_cnu_59_in_3, msg_to_check_it_1_cnu_85_in_3);
vnu variable_node_105_1(data_105, msg_to_bit_it_1_vnu_105_in_0, msg_to_bit_it_1_vnu_105_in_1, msg_to_bit_it_1_vnu_105_in_2, msg_to_check_it_1_cnu_30_in_3, msg_to_check_it_1_cnu_60_in_3, msg_to_check_it_1_cnu_86_in_3);
vnu variable_node_106_1(data_106, msg_to_bit_it_1_vnu_106_in_0, msg_to_bit_it_1_vnu_106_in_1, msg_to_bit_it_1_vnu_106_in_2, msg_to_check_it_1_cnu_31_in_3, msg_to_check_it_1_cnu_61_in_3, msg_to_check_it_1_cnu_87_in_3);
vnu variable_node_107_1(data_107, msg_to_bit_it_1_vnu_107_in_0, msg_to_bit_it_1_vnu_107_in_1, msg_to_bit_it_1_vnu_107_in_2, msg_to_check_it_1_cnu_32_in_3, msg_to_check_it_1_cnu_62_in_3, msg_to_check_it_1_cnu_88_in_3);
vnu variable_node_108_1(data_108, msg_to_bit_it_1_vnu_108_in_0, msg_to_bit_it_1_vnu_108_in_1, msg_to_bit_it_1_vnu_108_in_2, msg_to_check_it_1_cnu_0_in_3, msg_to_check_it_1_cnu_63_in_3, msg_to_check_it_1_cnu_89_in_3);
vnu variable_node_109_1(data_109, msg_to_bit_it_1_vnu_109_in_0, msg_to_bit_it_1_vnu_109_in_1, msg_to_bit_it_1_vnu_109_in_2, msg_to_check_it_1_cnu_1_in_3, msg_to_check_it_1_cnu_64_in_3, msg_to_check_it_1_cnu_90_in_3);
vnu variable_node_110_1(data_110, msg_to_bit_it_1_vnu_110_in_0, msg_to_bit_it_1_vnu_110_in_1, msg_to_bit_it_1_vnu_110_in_2, msg_to_check_it_1_cnu_2_in_3, msg_to_check_it_1_cnu_65_in_3, msg_to_check_it_1_cnu_91_in_3);
vnu variable_node_111_1(data_111, msg_to_bit_it_1_vnu_111_in_0, msg_to_bit_it_1_vnu_111_in_1, msg_to_bit_it_1_vnu_111_in_2, msg_to_check_it_1_cnu_3_in_3, msg_to_check_it_1_cnu_33_in_3, msg_to_check_it_1_cnu_92_in_3);
vnu variable_node_112_1(data_112, msg_to_bit_it_1_vnu_112_in_0, msg_to_bit_it_1_vnu_112_in_1, msg_to_bit_it_1_vnu_112_in_2, msg_to_check_it_1_cnu_4_in_3, msg_to_check_it_1_cnu_34_in_3, msg_to_check_it_1_cnu_93_in_3);
vnu variable_node_113_1(data_113, msg_to_bit_it_1_vnu_113_in_0, msg_to_bit_it_1_vnu_113_in_1, msg_to_bit_it_1_vnu_113_in_2, msg_to_check_it_1_cnu_5_in_3, msg_to_check_it_1_cnu_35_in_3, msg_to_check_it_1_cnu_94_in_3);
vnu variable_node_114_1(data_114, msg_to_bit_it_1_vnu_114_in_0, msg_to_bit_it_1_vnu_114_in_1, msg_to_bit_it_1_vnu_114_in_2, msg_to_check_it_1_cnu_6_in_3, msg_to_check_it_1_cnu_36_in_3, msg_to_check_it_1_cnu_95_in_3);
vnu variable_node_115_1(data_115, msg_to_bit_it_1_vnu_115_in_0, msg_to_bit_it_1_vnu_115_in_1, msg_to_bit_it_1_vnu_115_in_2, msg_to_check_it_1_cnu_7_in_3, msg_to_check_it_1_cnu_37_in_3, msg_to_check_it_1_cnu_96_in_3);
vnu variable_node_116_1(data_116, msg_to_bit_it_1_vnu_116_in_0, msg_to_bit_it_1_vnu_116_in_1, msg_to_bit_it_1_vnu_116_in_2, msg_to_check_it_1_cnu_8_in_3, msg_to_check_it_1_cnu_38_in_3, msg_to_check_it_1_cnu_97_in_3);
vnu variable_node_117_1(data_117, msg_to_bit_it_1_vnu_117_in_0, msg_to_bit_it_1_vnu_117_in_1, msg_to_bit_it_1_vnu_117_in_2, msg_to_check_it_1_cnu_9_in_3, msg_to_check_it_1_cnu_39_in_3, msg_to_check_it_1_cnu_98_in_3);
vnu variable_node_118_1(data_118, msg_to_bit_it_1_vnu_118_in_0, msg_to_bit_it_1_vnu_118_in_1, msg_to_bit_it_1_vnu_118_in_2, msg_to_check_it_1_cnu_10_in_3, msg_to_check_it_1_cnu_40_in_3, msg_to_check_it_1_cnu_66_in_3);
vnu variable_node_119_1(data_119, msg_to_bit_it_1_vnu_119_in_0, msg_to_bit_it_1_vnu_119_in_1, msg_to_bit_it_1_vnu_119_in_2, msg_to_check_it_1_cnu_11_in_3, msg_to_check_it_1_cnu_41_in_3, msg_to_check_it_1_cnu_67_in_3);
vnu variable_node_120_1(data_120, msg_to_bit_it_1_vnu_120_in_0, msg_to_bit_it_1_vnu_120_in_1, msg_to_bit_it_1_vnu_120_in_2, msg_to_check_it_1_cnu_12_in_3, msg_to_check_it_1_cnu_42_in_3, msg_to_check_it_1_cnu_68_in_3);
vnu variable_node_121_1(data_121, msg_to_bit_it_1_vnu_121_in_0, msg_to_bit_it_1_vnu_121_in_1, msg_to_bit_it_1_vnu_121_in_2, msg_to_check_it_1_cnu_13_in_3, msg_to_check_it_1_cnu_43_in_3, msg_to_check_it_1_cnu_69_in_3);
vnu variable_node_122_1(data_122, msg_to_bit_it_1_vnu_122_in_0, msg_to_bit_it_1_vnu_122_in_1, msg_to_bit_it_1_vnu_122_in_2, msg_to_check_it_1_cnu_14_in_3, msg_to_check_it_1_cnu_44_in_3, msg_to_check_it_1_cnu_70_in_3);
vnu variable_node_123_1(data_123, msg_to_bit_it_1_vnu_123_in_0, msg_to_bit_it_1_vnu_123_in_1, msg_to_bit_it_1_vnu_123_in_2, msg_to_check_it_1_cnu_15_in_3, msg_to_check_it_1_cnu_45_in_3, msg_to_check_it_1_cnu_71_in_3);
vnu variable_node_124_1(data_124, msg_to_bit_it_1_vnu_124_in_0, msg_to_bit_it_1_vnu_124_in_1, msg_to_bit_it_1_vnu_124_in_2, msg_to_check_it_1_cnu_16_in_3, msg_to_check_it_1_cnu_46_in_3, msg_to_check_it_1_cnu_72_in_3);
vnu variable_node_125_1(data_125, msg_to_bit_it_1_vnu_125_in_0, msg_to_bit_it_1_vnu_125_in_1, msg_to_bit_it_1_vnu_125_in_2, msg_to_check_it_1_cnu_17_in_3, msg_to_check_it_1_cnu_47_in_3, msg_to_check_it_1_cnu_73_in_3);
vnu variable_node_126_1(data_126, msg_to_bit_it_1_vnu_126_in_0, msg_to_bit_it_1_vnu_126_in_1, msg_to_bit_it_1_vnu_126_in_2, msg_to_check_it_1_cnu_18_in_3, msg_to_check_it_1_cnu_48_in_3, msg_to_check_it_1_cnu_74_in_3);
vnu variable_node_127_1(data_127, msg_to_bit_it_1_vnu_127_in_0, msg_to_bit_it_1_vnu_127_in_1, msg_to_bit_it_1_vnu_127_in_2, msg_to_check_it_1_cnu_19_in_3, msg_to_check_it_1_cnu_49_in_3, msg_to_check_it_1_cnu_75_in_3);
vnu variable_node_128_1(data_128, msg_to_bit_it_1_vnu_128_in_0, msg_to_bit_it_1_vnu_128_in_1, msg_to_bit_it_1_vnu_128_in_2, msg_to_check_it_1_cnu_20_in_3, msg_to_check_it_1_cnu_50_in_3, msg_to_check_it_1_cnu_76_in_3);
vnu variable_node_129_1(data_129, msg_to_bit_it_1_vnu_129_in_0, msg_to_bit_it_1_vnu_129_in_1, msg_to_bit_it_1_vnu_129_in_2, msg_to_check_it_1_cnu_21_in_3, msg_to_check_it_1_cnu_51_in_3, msg_to_check_it_1_cnu_77_in_3);
vnu variable_node_130_1(data_130, msg_to_bit_it_1_vnu_130_in_0, msg_to_bit_it_1_vnu_130_in_1, msg_to_bit_it_1_vnu_130_in_2, msg_to_check_it_1_cnu_22_in_3, msg_to_check_it_1_cnu_52_in_3, msg_to_check_it_1_cnu_78_in_3);
vnu variable_node_131_1(data_131, msg_to_bit_it_1_vnu_131_in_0, msg_to_bit_it_1_vnu_131_in_1, msg_to_bit_it_1_vnu_131_in_2, msg_to_check_it_1_cnu_23_in_3, msg_to_check_it_1_cnu_53_in_3, msg_to_check_it_1_cnu_79_in_3);
vnu variable_node_132_1(data_132, msg_to_bit_it_1_vnu_132_in_0, msg_to_bit_it_1_vnu_132_in_1, msg_to_bit_it_1_vnu_132_in_2, msg_to_check_it_1_cnu_18_in_4, msg_to_check_it_1_cnu_43_in_4, msg_to_check_it_1_cnu_72_in_4);
vnu variable_node_133_1(data_133, msg_to_bit_it_1_vnu_133_in_0, msg_to_bit_it_1_vnu_133_in_1, msg_to_bit_it_1_vnu_133_in_2, msg_to_check_it_1_cnu_19_in_4, msg_to_check_it_1_cnu_44_in_4, msg_to_check_it_1_cnu_73_in_4);
vnu variable_node_134_1(data_134, msg_to_bit_it_1_vnu_134_in_0, msg_to_bit_it_1_vnu_134_in_1, msg_to_bit_it_1_vnu_134_in_2, msg_to_check_it_1_cnu_20_in_4, msg_to_check_it_1_cnu_45_in_4, msg_to_check_it_1_cnu_74_in_4);
vnu variable_node_135_1(data_135, msg_to_bit_it_1_vnu_135_in_0, msg_to_bit_it_1_vnu_135_in_1, msg_to_bit_it_1_vnu_135_in_2, msg_to_check_it_1_cnu_21_in_4, msg_to_check_it_1_cnu_46_in_4, msg_to_check_it_1_cnu_75_in_4);
vnu variable_node_136_1(data_136, msg_to_bit_it_1_vnu_136_in_0, msg_to_bit_it_1_vnu_136_in_1, msg_to_bit_it_1_vnu_136_in_2, msg_to_check_it_1_cnu_22_in_4, msg_to_check_it_1_cnu_47_in_4, msg_to_check_it_1_cnu_76_in_4);
vnu variable_node_137_1(data_137, msg_to_bit_it_1_vnu_137_in_0, msg_to_bit_it_1_vnu_137_in_1, msg_to_bit_it_1_vnu_137_in_2, msg_to_check_it_1_cnu_23_in_4, msg_to_check_it_1_cnu_48_in_4, msg_to_check_it_1_cnu_77_in_4);
vnu variable_node_138_1(data_138, msg_to_bit_it_1_vnu_138_in_0, msg_to_bit_it_1_vnu_138_in_1, msg_to_bit_it_1_vnu_138_in_2, msg_to_check_it_1_cnu_24_in_4, msg_to_check_it_1_cnu_49_in_4, msg_to_check_it_1_cnu_78_in_4);
vnu variable_node_139_1(data_139, msg_to_bit_it_1_vnu_139_in_0, msg_to_bit_it_1_vnu_139_in_1, msg_to_bit_it_1_vnu_139_in_2, msg_to_check_it_1_cnu_25_in_4, msg_to_check_it_1_cnu_50_in_4, msg_to_check_it_1_cnu_79_in_4);
vnu variable_node_140_1(data_140, msg_to_bit_it_1_vnu_140_in_0, msg_to_bit_it_1_vnu_140_in_1, msg_to_bit_it_1_vnu_140_in_2, msg_to_check_it_1_cnu_26_in_4, msg_to_check_it_1_cnu_51_in_4, msg_to_check_it_1_cnu_80_in_4);
vnu variable_node_141_1(data_141, msg_to_bit_it_1_vnu_141_in_0, msg_to_bit_it_1_vnu_141_in_1, msg_to_bit_it_1_vnu_141_in_2, msg_to_check_it_1_cnu_27_in_4, msg_to_check_it_1_cnu_52_in_4, msg_to_check_it_1_cnu_81_in_4);
vnu variable_node_142_1(data_142, msg_to_bit_it_1_vnu_142_in_0, msg_to_bit_it_1_vnu_142_in_1, msg_to_bit_it_1_vnu_142_in_2, msg_to_check_it_1_cnu_28_in_4, msg_to_check_it_1_cnu_53_in_4, msg_to_check_it_1_cnu_82_in_4);
vnu variable_node_143_1(data_143, msg_to_bit_it_1_vnu_143_in_0, msg_to_bit_it_1_vnu_143_in_1, msg_to_bit_it_1_vnu_143_in_2, msg_to_check_it_1_cnu_29_in_4, msg_to_check_it_1_cnu_54_in_4, msg_to_check_it_1_cnu_83_in_4);
vnu variable_node_144_1(data_144, msg_to_bit_it_1_vnu_144_in_0, msg_to_bit_it_1_vnu_144_in_1, msg_to_bit_it_1_vnu_144_in_2, msg_to_check_it_1_cnu_30_in_4, msg_to_check_it_1_cnu_55_in_4, msg_to_check_it_1_cnu_84_in_4);
vnu variable_node_145_1(data_145, msg_to_bit_it_1_vnu_145_in_0, msg_to_bit_it_1_vnu_145_in_1, msg_to_bit_it_1_vnu_145_in_2, msg_to_check_it_1_cnu_31_in_4, msg_to_check_it_1_cnu_56_in_4, msg_to_check_it_1_cnu_85_in_4);
vnu variable_node_146_1(data_146, msg_to_bit_it_1_vnu_146_in_0, msg_to_bit_it_1_vnu_146_in_1, msg_to_bit_it_1_vnu_146_in_2, msg_to_check_it_1_cnu_32_in_4, msg_to_check_it_1_cnu_57_in_4, msg_to_check_it_1_cnu_86_in_4);
vnu variable_node_147_1(data_147, msg_to_bit_it_1_vnu_147_in_0, msg_to_bit_it_1_vnu_147_in_1, msg_to_bit_it_1_vnu_147_in_2, msg_to_check_it_1_cnu_0_in_4, msg_to_check_it_1_cnu_58_in_4, msg_to_check_it_1_cnu_87_in_4);
vnu variable_node_148_1(data_148, msg_to_bit_it_1_vnu_148_in_0, msg_to_bit_it_1_vnu_148_in_1, msg_to_bit_it_1_vnu_148_in_2, msg_to_check_it_1_cnu_1_in_4, msg_to_check_it_1_cnu_59_in_4, msg_to_check_it_1_cnu_88_in_4);
vnu variable_node_149_1(data_149, msg_to_bit_it_1_vnu_149_in_0, msg_to_bit_it_1_vnu_149_in_1, msg_to_bit_it_1_vnu_149_in_2, msg_to_check_it_1_cnu_2_in_4, msg_to_check_it_1_cnu_60_in_4, msg_to_check_it_1_cnu_89_in_4);
vnu variable_node_150_1(data_150, msg_to_bit_it_1_vnu_150_in_0, msg_to_bit_it_1_vnu_150_in_1, msg_to_bit_it_1_vnu_150_in_2, msg_to_check_it_1_cnu_3_in_4, msg_to_check_it_1_cnu_61_in_4, msg_to_check_it_1_cnu_90_in_4);
vnu variable_node_151_1(data_151, msg_to_bit_it_1_vnu_151_in_0, msg_to_bit_it_1_vnu_151_in_1, msg_to_bit_it_1_vnu_151_in_2, msg_to_check_it_1_cnu_4_in_4, msg_to_check_it_1_cnu_62_in_4, msg_to_check_it_1_cnu_91_in_4);
vnu variable_node_152_1(data_152, msg_to_bit_it_1_vnu_152_in_0, msg_to_bit_it_1_vnu_152_in_1, msg_to_bit_it_1_vnu_152_in_2, msg_to_check_it_1_cnu_5_in_4, msg_to_check_it_1_cnu_63_in_4, msg_to_check_it_1_cnu_92_in_4);
vnu variable_node_153_1(data_153, msg_to_bit_it_1_vnu_153_in_0, msg_to_bit_it_1_vnu_153_in_1, msg_to_bit_it_1_vnu_153_in_2, msg_to_check_it_1_cnu_6_in_4, msg_to_check_it_1_cnu_64_in_4, msg_to_check_it_1_cnu_93_in_4);
vnu variable_node_154_1(data_154, msg_to_bit_it_1_vnu_154_in_0, msg_to_bit_it_1_vnu_154_in_1, msg_to_bit_it_1_vnu_154_in_2, msg_to_check_it_1_cnu_7_in_4, msg_to_check_it_1_cnu_65_in_4, msg_to_check_it_1_cnu_94_in_4);
vnu variable_node_155_1(data_155, msg_to_bit_it_1_vnu_155_in_0, msg_to_bit_it_1_vnu_155_in_1, msg_to_bit_it_1_vnu_155_in_2, msg_to_check_it_1_cnu_8_in_4, msg_to_check_it_1_cnu_33_in_4, msg_to_check_it_1_cnu_95_in_4);
vnu variable_node_156_1(data_156, msg_to_bit_it_1_vnu_156_in_0, msg_to_bit_it_1_vnu_156_in_1, msg_to_bit_it_1_vnu_156_in_2, msg_to_check_it_1_cnu_9_in_4, msg_to_check_it_1_cnu_34_in_4, msg_to_check_it_1_cnu_96_in_4);
vnu variable_node_157_1(data_157, msg_to_bit_it_1_vnu_157_in_0, msg_to_bit_it_1_vnu_157_in_1, msg_to_bit_it_1_vnu_157_in_2, msg_to_check_it_1_cnu_10_in_4, msg_to_check_it_1_cnu_35_in_4, msg_to_check_it_1_cnu_97_in_4);
vnu variable_node_158_1(data_158, msg_to_bit_it_1_vnu_158_in_0, msg_to_bit_it_1_vnu_158_in_1, msg_to_bit_it_1_vnu_158_in_2, msg_to_check_it_1_cnu_11_in_4, msg_to_check_it_1_cnu_36_in_4, msg_to_check_it_1_cnu_98_in_4);
vnu variable_node_159_1(data_159, msg_to_bit_it_1_vnu_159_in_0, msg_to_bit_it_1_vnu_159_in_1, msg_to_bit_it_1_vnu_159_in_2, msg_to_check_it_1_cnu_12_in_4, msg_to_check_it_1_cnu_37_in_4, msg_to_check_it_1_cnu_66_in_4);
vnu variable_node_160_1(data_160, msg_to_bit_it_1_vnu_160_in_0, msg_to_bit_it_1_vnu_160_in_1, msg_to_bit_it_1_vnu_160_in_2, msg_to_check_it_1_cnu_13_in_4, msg_to_check_it_1_cnu_38_in_4, msg_to_check_it_1_cnu_67_in_4);
vnu variable_node_161_1(data_161, msg_to_bit_it_1_vnu_161_in_0, msg_to_bit_it_1_vnu_161_in_1, msg_to_bit_it_1_vnu_161_in_2, msg_to_check_it_1_cnu_14_in_4, msg_to_check_it_1_cnu_39_in_4, msg_to_check_it_1_cnu_68_in_4);
vnu variable_node_162_1(data_162, msg_to_bit_it_1_vnu_162_in_0, msg_to_bit_it_1_vnu_162_in_1, msg_to_bit_it_1_vnu_162_in_2, msg_to_check_it_1_cnu_15_in_4, msg_to_check_it_1_cnu_40_in_4, msg_to_check_it_1_cnu_69_in_4);
vnu variable_node_163_1(data_163, msg_to_bit_it_1_vnu_163_in_0, msg_to_bit_it_1_vnu_163_in_1, msg_to_bit_it_1_vnu_163_in_2, msg_to_check_it_1_cnu_16_in_4, msg_to_check_it_1_cnu_41_in_4, msg_to_check_it_1_cnu_70_in_4);
vnu variable_node_164_1(data_164, msg_to_bit_it_1_vnu_164_in_0, msg_to_bit_it_1_vnu_164_in_1, msg_to_bit_it_1_vnu_164_in_2, msg_to_check_it_1_cnu_17_in_4, msg_to_check_it_1_cnu_42_in_4, msg_to_check_it_1_cnu_71_in_4);
vnu variable_node_165_1(data_165, msg_to_bit_it_1_vnu_165_in_0, msg_to_bit_it_1_vnu_165_in_1, msg_to_bit_it_1_vnu_165_in_2, msg_to_check_it_1_cnu_13_in_5, msg_to_check_it_1_cnu_41_in_5, msg_to_check_it_1_cnu_69_in_5);
vnu variable_node_166_1(data_166, msg_to_bit_it_1_vnu_166_in_0, msg_to_bit_it_1_vnu_166_in_1, msg_to_bit_it_1_vnu_166_in_2, msg_to_check_it_1_cnu_14_in_5, msg_to_check_it_1_cnu_42_in_5, msg_to_check_it_1_cnu_70_in_5);
vnu variable_node_167_1(data_167, msg_to_bit_it_1_vnu_167_in_0, msg_to_bit_it_1_vnu_167_in_1, msg_to_bit_it_1_vnu_167_in_2, msg_to_check_it_1_cnu_15_in_5, msg_to_check_it_1_cnu_43_in_5, msg_to_check_it_1_cnu_71_in_5);
vnu variable_node_168_1(data_168, msg_to_bit_it_1_vnu_168_in_0, msg_to_bit_it_1_vnu_168_in_1, msg_to_bit_it_1_vnu_168_in_2, msg_to_check_it_1_cnu_16_in_5, msg_to_check_it_1_cnu_44_in_5, msg_to_check_it_1_cnu_72_in_5);
vnu variable_node_169_1(data_169, msg_to_bit_it_1_vnu_169_in_0, msg_to_bit_it_1_vnu_169_in_1, msg_to_bit_it_1_vnu_169_in_2, msg_to_check_it_1_cnu_17_in_5, msg_to_check_it_1_cnu_45_in_5, msg_to_check_it_1_cnu_73_in_5);
vnu variable_node_170_1(data_170, msg_to_bit_it_1_vnu_170_in_0, msg_to_bit_it_1_vnu_170_in_1, msg_to_bit_it_1_vnu_170_in_2, msg_to_check_it_1_cnu_18_in_5, msg_to_check_it_1_cnu_46_in_5, msg_to_check_it_1_cnu_74_in_5);
vnu variable_node_171_1(data_171, msg_to_bit_it_1_vnu_171_in_0, msg_to_bit_it_1_vnu_171_in_1, msg_to_bit_it_1_vnu_171_in_2, msg_to_check_it_1_cnu_19_in_5, msg_to_check_it_1_cnu_47_in_5, msg_to_check_it_1_cnu_75_in_5);
vnu variable_node_172_1(data_172, msg_to_bit_it_1_vnu_172_in_0, msg_to_bit_it_1_vnu_172_in_1, msg_to_bit_it_1_vnu_172_in_2, msg_to_check_it_1_cnu_20_in_5, msg_to_check_it_1_cnu_48_in_5, msg_to_check_it_1_cnu_76_in_5);
vnu variable_node_173_1(data_173, msg_to_bit_it_1_vnu_173_in_0, msg_to_bit_it_1_vnu_173_in_1, msg_to_bit_it_1_vnu_173_in_2, msg_to_check_it_1_cnu_21_in_5, msg_to_check_it_1_cnu_49_in_5, msg_to_check_it_1_cnu_77_in_5);
vnu variable_node_174_1(data_174, msg_to_bit_it_1_vnu_174_in_0, msg_to_bit_it_1_vnu_174_in_1, msg_to_bit_it_1_vnu_174_in_2, msg_to_check_it_1_cnu_22_in_5, msg_to_check_it_1_cnu_50_in_5, msg_to_check_it_1_cnu_78_in_5);
vnu variable_node_175_1(data_175, msg_to_bit_it_1_vnu_175_in_0, msg_to_bit_it_1_vnu_175_in_1, msg_to_bit_it_1_vnu_175_in_2, msg_to_check_it_1_cnu_23_in_5, msg_to_check_it_1_cnu_51_in_5, msg_to_check_it_1_cnu_79_in_5);
vnu variable_node_176_1(data_176, msg_to_bit_it_1_vnu_176_in_0, msg_to_bit_it_1_vnu_176_in_1, msg_to_bit_it_1_vnu_176_in_2, msg_to_check_it_1_cnu_24_in_5, msg_to_check_it_1_cnu_52_in_5, msg_to_check_it_1_cnu_80_in_5);
vnu variable_node_177_1(data_177, msg_to_bit_it_1_vnu_177_in_0, msg_to_bit_it_1_vnu_177_in_1, msg_to_bit_it_1_vnu_177_in_2, msg_to_check_it_1_cnu_25_in_5, msg_to_check_it_1_cnu_53_in_5, msg_to_check_it_1_cnu_81_in_5);
vnu variable_node_178_1(data_178, msg_to_bit_it_1_vnu_178_in_0, msg_to_bit_it_1_vnu_178_in_1, msg_to_bit_it_1_vnu_178_in_2, msg_to_check_it_1_cnu_26_in_5, msg_to_check_it_1_cnu_54_in_5, msg_to_check_it_1_cnu_82_in_5);
vnu variable_node_179_1(data_179, msg_to_bit_it_1_vnu_179_in_0, msg_to_bit_it_1_vnu_179_in_1, msg_to_bit_it_1_vnu_179_in_2, msg_to_check_it_1_cnu_27_in_5, msg_to_check_it_1_cnu_55_in_5, msg_to_check_it_1_cnu_83_in_5);
vnu variable_node_180_1(data_180, msg_to_bit_it_1_vnu_180_in_0, msg_to_bit_it_1_vnu_180_in_1, msg_to_bit_it_1_vnu_180_in_2, msg_to_check_it_1_cnu_28_in_5, msg_to_check_it_1_cnu_56_in_5, msg_to_check_it_1_cnu_84_in_5);
vnu variable_node_181_1(data_181, msg_to_bit_it_1_vnu_181_in_0, msg_to_bit_it_1_vnu_181_in_1, msg_to_bit_it_1_vnu_181_in_2, msg_to_check_it_1_cnu_29_in_5, msg_to_check_it_1_cnu_57_in_5, msg_to_check_it_1_cnu_85_in_5);
vnu variable_node_182_1(data_182, msg_to_bit_it_1_vnu_182_in_0, msg_to_bit_it_1_vnu_182_in_1, msg_to_bit_it_1_vnu_182_in_2, msg_to_check_it_1_cnu_30_in_5, msg_to_check_it_1_cnu_58_in_5, msg_to_check_it_1_cnu_86_in_5);
vnu variable_node_183_1(data_183, msg_to_bit_it_1_vnu_183_in_0, msg_to_bit_it_1_vnu_183_in_1, msg_to_bit_it_1_vnu_183_in_2, msg_to_check_it_1_cnu_31_in_5, msg_to_check_it_1_cnu_59_in_5, msg_to_check_it_1_cnu_87_in_5);
vnu variable_node_184_1(data_184, msg_to_bit_it_1_vnu_184_in_0, msg_to_bit_it_1_vnu_184_in_1, msg_to_bit_it_1_vnu_184_in_2, msg_to_check_it_1_cnu_32_in_5, msg_to_check_it_1_cnu_60_in_5, msg_to_check_it_1_cnu_88_in_5);
vnu variable_node_185_1(data_185, msg_to_bit_it_1_vnu_185_in_0, msg_to_bit_it_1_vnu_185_in_1, msg_to_bit_it_1_vnu_185_in_2, msg_to_check_it_1_cnu_0_in_5, msg_to_check_it_1_cnu_61_in_5, msg_to_check_it_1_cnu_89_in_5);
vnu variable_node_186_1(data_186, msg_to_bit_it_1_vnu_186_in_0, msg_to_bit_it_1_vnu_186_in_1, msg_to_bit_it_1_vnu_186_in_2, msg_to_check_it_1_cnu_1_in_5, msg_to_check_it_1_cnu_62_in_5, msg_to_check_it_1_cnu_90_in_5);
vnu variable_node_187_1(data_187, msg_to_bit_it_1_vnu_187_in_0, msg_to_bit_it_1_vnu_187_in_1, msg_to_bit_it_1_vnu_187_in_2, msg_to_check_it_1_cnu_2_in_5, msg_to_check_it_1_cnu_63_in_5, msg_to_check_it_1_cnu_91_in_5);
vnu variable_node_188_1(data_188, msg_to_bit_it_1_vnu_188_in_0, msg_to_bit_it_1_vnu_188_in_1, msg_to_bit_it_1_vnu_188_in_2, msg_to_check_it_1_cnu_3_in_5, msg_to_check_it_1_cnu_64_in_5, msg_to_check_it_1_cnu_92_in_5);
vnu variable_node_189_1(data_189, msg_to_bit_it_1_vnu_189_in_0, msg_to_bit_it_1_vnu_189_in_1, msg_to_bit_it_1_vnu_189_in_2, msg_to_check_it_1_cnu_4_in_5, msg_to_check_it_1_cnu_65_in_5, msg_to_check_it_1_cnu_93_in_5);
vnu variable_node_190_1(data_190, msg_to_bit_it_1_vnu_190_in_0, msg_to_bit_it_1_vnu_190_in_1, msg_to_bit_it_1_vnu_190_in_2, msg_to_check_it_1_cnu_5_in_5, msg_to_check_it_1_cnu_33_in_5, msg_to_check_it_1_cnu_94_in_5);
vnu variable_node_191_1(data_191, msg_to_bit_it_1_vnu_191_in_0, msg_to_bit_it_1_vnu_191_in_1, msg_to_bit_it_1_vnu_191_in_2, msg_to_check_it_1_cnu_6_in_5, msg_to_check_it_1_cnu_34_in_5, msg_to_check_it_1_cnu_95_in_5);
vnu variable_node_192_1(data_192, msg_to_bit_it_1_vnu_192_in_0, msg_to_bit_it_1_vnu_192_in_1, msg_to_bit_it_1_vnu_192_in_2, msg_to_check_it_1_cnu_7_in_5, msg_to_check_it_1_cnu_35_in_5, msg_to_check_it_1_cnu_96_in_5);
vnu variable_node_193_1(data_193, msg_to_bit_it_1_vnu_193_in_0, msg_to_bit_it_1_vnu_193_in_1, msg_to_bit_it_1_vnu_193_in_2, msg_to_check_it_1_cnu_8_in_5, msg_to_check_it_1_cnu_36_in_5, msg_to_check_it_1_cnu_97_in_5);
vnu variable_node_194_1(data_194, msg_to_bit_it_1_vnu_194_in_0, msg_to_bit_it_1_vnu_194_in_1, msg_to_bit_it_1_vnu_194_in_2, msg_to_check_it_1_cnu_9_in_5, msg_to_check_it_1_cnu_37_in_5, msg_to_check_it_1_cnu_98_in_5);
vnu variable_node_195_1(data_195, msg_to_bit_it_1_vnu_195_in_0, msg_to_bit_it_1_vnu_195_in_1, msg_to_bit_it_1_vnu_195_in_2, msg_to_check_it_1_cnu_10_in_5, msg_to_check_it_1_cnu_38_in_5, msg_to_check_it_1_cnu_66_in_5);
vnu variable_node_196_1(data_196, msg_to_bit_it_1_vnu_196_in_0, msg_to_bit_it_1_vnu_196_in_1, msg_to_bit_it_1_vnu_196_in_2, msg_to_check_it_1_cnu_11_in_5, msg_to_check_it_1_cnu_39_in_5, msg_to_check_it_1_cnu_67_in_5);
vnu variable_node_197_1(data_197, msg_to_bit_it_1_vnu_197_in_0, msg_to_bit_it_1_vnu_197_in_1, msg_to_bit_it_1_vnu_197_in_2, msg_to_check_it_1_cnu_12_in_5, msg_to_check_it_1_cnu_40_in_5, msg_to_check_it_1_cnu_68_in_5);



cnu check_node_0_1(msg_to_check_it_1_cnu_0_in_0, msg_to_check_it_1_cnu_0_in_1, msg_to_check_it_1_cnu_0_in_2, msg_to_check_it_1_cnu_0_in_3, msg_to_check_it_1_cnu_0_in_4, msg_to_check_it_1_cnu_0_in_5, msg_to_bit_it_2_vnu_2_in_0, msg_to_bit_it_2_vnu_36_in_0, msg_to_bit_it_2_vnu_73_in_0, msg_to_bit_it_2_vnu_108_in_0, msg_to_bit_it_2_vnu_147_in_0, msg_to_bit_it_2_vnu_185_in_0);
cnu check_node_1_1(msg_to_check_it_1_cnu_1_in_0, msg_to_check_it_1_cnu_1_in_1, msg_to_check_it_1_cnu_1_in_2, msg_to_check_it_1_cnu_1_in_3, msg_to_check_it_1_cnu_1_in_4, msg_to_check_it_1_cnu_1_in_5, msg_to_bit_it_2_vnu_3_in_0, msg_to_bit_it_2_vnu_37_in_0, msg_to_bit_it_2_vnu_74_in_0, msg_to_bit_it_2_vnu_109_in_0, msg_to_bit_it_2_vnu_148_in_0, msg_to_bit_it_2_vnu_186_in_0);
cnu check_node_2_1(msg_to_check_it_1_cnu_2_in_0, msg_to_check_it_1_cnu_2_in_1, msg_to_check_it_1_cnu_2_in_2, msg_to_check_it_1_cnu_2_in_3, msg_to_check_it_1_cnu_2_in_4, msg_to_check_it_1_cnu_2_in_5, msg_to_bit_it_2_vnu_4_in_0, msg_to_bit_it_2_vnu_38_in_0, msg_to_bit_it_2_vnu_75_in_0, msg_to_bit_it_2_vnu_110_in_0, msg_to_bit_it_2_vnu_149_in_0, msg_to_bit_it_2_vnu_187_in_0);
cnu check_node_3_1(msg_to_check_it_1_cnu_3_in_0, msg_to_check_it_1_cnu_3_in_1, msg_to_check_it_1_cnu_3_in_2, msg_to_check_it_1_cnu_3_in_3, msg_to_check_it_1_cnu_3_in_4, msg_to_check_it_1_cnu_3_in_5, msg_to_bit_it_2_vnu_5_in_0, msg_to_bit_it_2_vnu_39_in_0, msg_to_bit_it_2_vnu_76_in_0, msg_to_bit_it_2_vnu_111_in_0, msg_to_bit_it_2_vnu_150_in_0, msg_to_bit_it_2_vnu_188_in_0);
cnu check_node_4_1(msg_to_check_it_1_cnu_4_in_0, msg_to_check_it_1_cnu_4_in_1, msg_to_check_it_1_cnu_4_in_2, msg_to_check_it_1_cnu_4_in_3, msg_to_check_it_1_cnu_4_in_4, msg_to_check_it_1_cnu_4_in_5, msg_to_bit_it_2_vnu_6_in_0, msg_to_bit_it_2_vnu_40_in_0, msg_to_bit_it_2_vnu_77_in_0, msg_to_bit_it_2_vnu_112_in_0, msg_to_bit_it_2_vnu_151_in_0, msg_to_bit_it_2_vnu_189_in_0);
cnu check_node_5_1(msg_to_check_it_1_cnu_5_in_0, msg_to_check_it_1_cnu_5_in_1, msg_to_check_it_1_cnu_5_in_2, msg_to_check_it_1_cnu_5_in_3, msg_to_check_it_1_cnu_5_in_4, msg_to_check_it_1_cnu_5_in_5, msg_to_bit_it_2_vnu_7_in_0, msg_to_bit_it_2_vnu_41_in_0, msg_to_bit_it_2_vnu_78_in_0, msg_to_bit_it_2_vnu_113_in_0, msg_to_bit_it_2_vnu_152_in_0, msg_to_bit_it_2_vnu_190_in_0);
cnu check_node_6_1(msg_to_check_it_1_cnu_6_in_0, msg_to_check_it_1_cnu_6_in_1, msg_to_check_it_1_cnu_6_in_2, msg_to_check_it_1_cnu_6_in_3, msg_to_check_it_1_cnu_6_in_4, msg_to_check_it_1_cnu_6_in_5, msg_to_bit_it_2_vnu_8_in_0, msg_to_bit_it_2_vnu_42_in_0, msg_to_bit_it_2_vnu_79_in_0, msg_to_bit_it_2_vnu_114_in_0, msg_to_bit_it_2_vnu_153_in_0, msg_to_bit_it_2_vnu_191_in_0);
cnu check_node_7_1(msg_to_check_it_1_cnu_7_in_0, msg_to_check_it_1_cnu_7_in_1, msg_to_check_it_1_cnu_7_in_2, msg_to_check_it_1_cnu_7_in_3, msg_to_check_it_1_cnu_7_in_4, msg_to_check_it_1_cnu_7_in_5, msg_to_bit_it_2_vnu_9_in_0, msg_to_bit_it_2_vnu_43_in_0, msg_to_bit_it_2_vnu_80_in_0, msg_to_bit_it_2_vnu_115_in_0, msg_to_bit_it_2_vnu_154_in_0, msg_to_bit_it_2_vnu_192_in_0);
cnu check_node_8_1(msg_to_check_it_1_cnu_8_in_0, msg_to_check_it_1_cnu_8_in_1, msg_to_check_it_1_cnu_8_in_2, msg_to_check_it_1_cnu_8_in_3, msg_to_check_it_1_cnu_8_in_4, msg_to_check_it_1_cnu_8_in_5, msg_to_bit_it_2_vnu_10_in_0, msg_to_bit_it_2_vnu_44_in_0, msg_to_bit_it_2_vnu_81_in_0, msg_to_bit_it_2_vnu_116_in_0, msg_to_bit_it_2_vnu_155_in_0, msg_to_bit_it_2_vnu_193_in_0);
cnu check_node_9_1(msg_to_check_it_1_cnu_9_in_0, msg_to_check_it_1_cnu_9_in_1, msg_to_check_it_1_cnu_9_in_2, msg_to_check_it_1_cnu_9_in_3, msg_to_check_it_1_cnu_9_in_4, msg_to_check_it_1_cnu_9_in_5, msg_to_bit_it_2_vnu_11_in_0, msg_to_bit_it_2_vnu_45_in_0, msg_to_bit_it_2_vnu_82_in_0, msg_to_bit_it_2_vnu_117_in_0, msg_to_bit_it_2_vnu_156_in_0, msg_to_bit_it_2_vnu_194_in_0);
cnu check_node_10_1(msg_to_check_it_1_cnu_10_in_0, msg_to_check_it_1_cnu_10_in_1, msg_to_check_it_1_cnu_10_in_2, msg_to_check_it_1_cnu_10_in_3, msg_to_check_it_1_cnu_10_in_4, msg_to_check_it_1_cnu_10_in_5, msg_to_bit_it_2_vnu_12_in_0, msg_to_bit_it_2_vnu_46_in_0, msg_to_bit_it_2_vnu_83_in_0, msg_to_bit_it_2_vnu_118_in_0, msg_to_bit_it_2_vnu_157_in_0, msg_to_bit_it_2_vnu_195_in_0);
cnu check_node_11_1(msg_to_check_it_1_cnu_11_in_0, msg_to_check_it_1_cnu_11_in_1, msg_to_check_it_1_cnu_11_in_2, msg_to_check_it_1_cnu_11_in_3, msg_to_check_it_1_cnu_11_in_4, msg_to_check_it_1_cnu_11_in_5, msg_to_bit_it_2_vnu_13_in_0, msg_to_bit_it_2_vnu_47_in_0, msg_to_bit_it_2_vnu_84_in_0, msg_to_bit_it_2_vnu_119_in_0, msg_to_bit_it_2_vnu_158_in_0, msg_to_bit_it_2_vnu_196_in_0);
cnu check_node_12_1(msg_to_check_it_1_cnu_12_in_0, msg_to_check_it_1_cnu_12_in_1, msg_to_check_it_1_cnu_12_in_2, msg_to_check_it_1_cnu_12_in_3, msg_to_check_it_1_cnu_12_in_4, msg_to_check_it_1_cnu_12_in_5, msg_to_bit_it_2_vnu_14_in_0, msg_to_bit_it_2_vnu_48_in_0, msg_to_bit_it_2_vnu_85_in_0, msg_to_bit_it_2_vnu_120_in_0, msg_to_bit_it_2_vnu_159_in_0, msg_to_bit_it_2_vnu_197_in_0);
cnu check_node_13_1(msg_to_check_it_1_cnu_13_in_0, msg_to_check_it_1_cnu_13_in_1, msg_to_check_it_1_cnu_13_in_2, msg_to_check_it_1_cnu_13_in_3, msg_to_check_it_1_cnu_13_in_4, msg_to_check_it_1_cnu_13_in_5, msg_to_bit_it_2_vnu_15_in_0, msg_to_bit_it_2_vnu_49_in_0, msg_to_bit_it_2_vnu_86_in_0, msg_to_bit_it_2_vnu_121_in_0, msg_to_bit_it_2_vnu_160_in_0, msg_to_bit_it_2_vnu_165_in_0);
cnu check_node_14_1(msg_to_check_it_1_cnu_14_in_0, msg_to_check_it_1_cnu_14_in_1, msg_to_check_it_1_cnu_14_in_2, msg_to_check_it_1_cnu_14_in_3, msg_to_check_it_1_cnu_14_in_4, msg_to_check_it_1_cnu_14_in_5, msg_to_bit_it_2_vnu_16_in_0, msg_to_bit_it_2_vnu_50_in_0, msg_to_bit_it_2_vnu_87_in_0, msg_to_bit_it_2_vnu_122_in_0, msg_to_bit_it_2_vnu_161_in_0, msg_to_bit_it_2_vnu_166_in_0);
cnu check_node_15_1(msg_to_check_it_1_cnu_15_in_0, msg_to_check_it_1_cnu_15_in_1, msg_to_check_it_1_cnu_15_in_2, msg_to_check_it_1_cnu_15_in_3, msg_to_check_it_1_cnu_15_in_4, msg_to_check_it_1_cnu_15_in_5, msg_to_bit_it_2_vnu_17_in_0, msg_to_bit_it_2_vnu_51_in_0, msg_to_bit_it_2_vnu_88_in_0, msg_to_bit_it_2_vnu_123_in_0, msg_to_bit_it_2_vnu_162_in_0, msg_to_bit_it_2_vnu_167_in_0);
cnu check_node_16_1(msg_to_check_it_1_cnu_16_in_0, msg_to_check_it_1_cnu_16_in_1, msg_to_check_it_1_cnu_16_in_2, msg_to_check_it_1_cnu_16_in_3, msg_to_check_it_1_cnu_16_in_4, msg_to_check_it_1_cnu_16_in_5, msg_to_bit_it_2_vnu_18_in_0, msg_to_bit_it_2_vnu_52_in_0, msg_to_bit_it_2_vnu_89_in_0, msg_to_bit_it_2_vnu_124_in_0, msg_to_bit_it_2_vnu_163_in_0, msg_to_bit_it_2_vnu_168_in_0);
cnu check_node_17_1(msg_to_check_it_1_cnu_17_in_0, msg_to_check_it_1_cnu_17_in_1, msg_to_check_it_1_cnu_17_in_2, msg_to_check_it_1_cnu_17_in_3, msg_to_check_it_1_cnu_17_in_4, msg_to_check_it_1_cnu_17_in_5, msg_to_bit_it_2_vnu_19_in_0, msg_to_bit_it_2_vnu_53_in_0, msg_to_bit_it_2_vnu_90_in_0, msg_to_bit_it_2_vnu_125_in_0, msg_to_bit_it_2_vnu_164_in_0, msg_to_bit_it_2_vnu_169_in_0);
cnu check_node_18_1(msg_to_check_it_1_cnu_18_in_0, msg_to_check_it_1_cnu_18_in_1, msg_to_check_it_1_cnu_18_in_2, msg_to_check_it_1_cnu_18_in_3, msg_to_check_it_1_cnu_18_in_4, msg_to_check_it_1_cnu_18_in_5, msg_to_bit_it_2_vnu_20_in_0, msg_to_bit_it_2_vnu_54_in_0, msg_to_bit_it_2_vnu_91_in_0, msg_to_bit_it_2_vnu_126_in_0, msg_to_bit_it_2_vnu_132_in_0, msg_to_bit_it_2_vnu_170_in_0);
cnu check_node_19_1(msg_to_check_it_1_cnu_19_in_0, msg_to_check_it_1_cnu_19_in_1, msg_to_check_it_1_cnu_19_in_2, msg_to_check_it_1_cnu_19_in_3, msg_to_check_it_1_cnu_19_in_4, msg_to_check_it_1_cnu_19_in_5, msg_to_bit_it_2_vnu_21_in_0, msg_to_bit_it_2_vnu_55_in_0, msg_to_bit_it_2_vnu_92_in_0, msg_to_bit_it_2_vnu_127_in_0, msg_to_bit_it_2_vnu_133_in_0, msg_to_bit_it_2_vnu_171_in_0);
cnu check_node_20_1(msg_to_check_it_1_cnu_20_in_0, msg_to_check_it_1_cnu_20_in_1, msg_to_check_it_1_cnu_20_in_2, msg_to_check_it_1_cnu_20_in_3, msg_to_check_it_1_cnu_20_in_4, msg_to_check_it_1_cnu_20_in_5, msg_to_bit_it_2_vnu_22_in_0, msg_to_bit_it_2_vnu_56_in_0, msg_to_bit_it_2_vnu_93_in_0, msg_to_bit_it_2_vnu_128_in_0, msg_to_bit_it_2_vnu_134_in_0, msg_to_bit_it_2_vnu_172_in_0);
cnu check_node_21_1(msg_to_check_it_1_cnu_21_in_0, msg_to_check_it_1_cnu_21_in_1, msg_to_check_it_1_cnu_21_in_2, msg_to_check_it_1_cnu_21_in_3, msg_to_check_it_1_cnu_21_in_4, msg_to_check_it_1_cnu_21_in_5, msg_to_bit_it_2_vnu_23_in_0, msg_to_bit_it_2_vnu_57_in_0, msg_to_bit_it_2_vnu_94_in_0, msg_to_bit_it_2_vnu_129_in_0, msg_to_bit_it_2_vnu_135_in_0, msg_to_bit_it_2_vnu_173_in_0);
cnu check_node_22_1(msg_to_check_it_1_cnu_22_in_0, msg_to_check_it_1_cnu_22_in_1, msg_to_check_it_1_cnu_22_in_2, msg_to_check_it_1_cnu_22_in_3, msg_to_check_it_1_cnu_22_in_4, msg_to_check_it_1_cnu_22_in_5, msg_to_bit_it_2_vnu_24_in_0, msg_to_bit_it_2_vnu_58_in_0, msg_to_bit_it_2_vnu_95_in_0, msg_to_bit_it_2_vnu_130_in_0, msg_to_bit_it_2_vnu_136_in_0, msg_to_bit_it_2_vnu_174_in_0);
cnu check_node_23_1(msg_to_check_it_1_cnu_23_in_0, msg_to_check_it_1_cnu_23_in_1, msg_to_check_it_1_cnu_23_in_2, msg_to_check_it_1_cnu_23_in_3, msg_to_check_it_1_cnu_23_in_4, msg_to_check_it_1_cnu_23_in_5, msg_to_bit_it_2_vnu_25_in_0, msg_to_bit_it_2_vnu_59_in_0, msg_to_bit_it_2_vnu_96_in_0, msg_to_bit_it_2_vnu_131_in_0, msg_to_bit_it_2_vnu_137_in_0, msg_to_bit_it_2_vnu_175_in_0);
cnu check_node_24_1(msg_to_check_it_1_cnu_24_in_0, msg_to_check_it_1_cnu_24_in_1, msg_to_check_it_1_cnu_24_in_2, msg_to_check_it_1_cnu_24_in_3, msg_to_check_it_1_cnu_24_in_4, msg_to_check_it_1_cnu_24_in_5, msg_to_bit_it_2_vnu_26_in_0, msg_to_bit_it_2_vnu_60_in_0, msg_to_bit_it_2_vnu_97_in_0, msg_to_bit_it_2_vnu_99_in_0, msg_to_bit_it_2_vnu_138_in_0, msg_to_bit_it_2_vnu_176_in_0);
cnu check_node_25_1(msg_to_check_it_1_cnu_25_in_0, msg_to_check_it_1_cnu_25_in_1, msg_to_check_it_1_cnu_25_in_2, msg_to_check_it_1_cnu_25_in_3, msg_to_check_it_1_cnu_25_in_4, msg_to_check_it_1_cnu_25_in_5, msg_to_bit_it_2_vnu_27_in_0, msg_to_bit_it_2_vnu_61_in_0, msg_to_bit_it_2_vnu_98_in_0, msg_to_bit_it_2_vnu_100_in_0, msg_to_bit_it_2_vnu_139_in_0, msg_to_bit_it_2_vnu_177_in_0);
cnu check_node_26_1(msg_to_check_it_1_cnu_26_in_0, msg_to_check_it_1_cnu_26_in_1, msg_to_check_it_1_cnu_26_in_2, msg_to_check_it_1_cnu_26_in_3, msg_to_check_it_1_cnu_26_in_4, msg_to_check_it_1_cnu_26_in_5, msg_to_bit_it_2_vnu_28_in_0, msg_to_bit_it_2_vnu_62_in_0, msg_to_bit_it_2_vnu_66_in_0, msg_to_bit_it_2_vnu_101_in_0, msg_to_bit_it_2_vnu_140_in_0, msg_to_bit_it_2_vnu_178_in_0);
cnu check_node_27_1(msg_to_check_it_1_cnu_27_in_0, msg_to_check_it_1_cnu_27_in_1, msg_to_check_it_1_cnu_27_in_2, msg_to_check_it_1_cnu_27_in_3, msg_to_check_it_1_cnu_27_in_4, msg_to_check_it_1_cnu_27_in_5, msg_to_bit_it_2_vnu_29_in_0, msg_to_bit_it_2_vnu_63_in_0, msg_to_bit_it_2_vnu_67_in_0, msg_to_bit_it_2_vnu_102_in_0, msg_to_bit_it_2_vnu_141_in_0, msg_to_bit_it_2_vnu_179_in_0);
cnu check_node_28_1(msg_to_check_it_1_cnu_28_in_0, msg_to_check_it_1_cnu_28_in_1, msg_to_check_it_1_cnu_28_in_2, msg_to_check_it_1_cnu_28_in_3, msg_to_check_it_1_cnu_28_in_4, msg_to_check_it_1_cnu_28_in_5, msg_to_bit_it_2_vnu_30_in_0, msg_to_bit_it_2_vnu_64_in_0, msg_to_bit_it_2_vnu_68_in_0, msg_to_bit_it_2_vnu_103_in_0, msg_to_bit_it_2_vnu_142_in_0, msg_to_bit_it_2_vnu_180_in_0);
cnu check_node_29_1(msg_to_check_it_1_cnu_29_in_0, msg_to_check_it_1_cnu_29_in_1, msg_to_check_it_1_cnu_29_in_2, msg_to_check_it_1_cnu_29_in_3, msg_to_check_it_1_cnu_29_in_4, msg_to_check_it_1_cnu_29_in_5, msg_to_bit_it_2_vnu_31_in_0, msg_to_bit_it_2_vnu_65_in_0, msg_to_bit_it_2_vnu_69_in_0, msg_to_bit_it_2_vnu_104_in_0, msg_to_bit_it_2_vnu_143_in_0, msg_to_bit_it_2_vnu_181_in_0);
cnu check_node_30_1(msg_to_check_it_1_cnu_30_in_0, msg_to_check_it_1_cnu_30_in_1, msg_to_check_it_1_cnu_30_in_2, msg_to_check_it_1_cnu_30_in_3, msg_to_check_it_1_cnu_30_in_4, msg_to_check_it_1_cnu_30_in_5, msg_to_bit_it_2_vnu_32_in_0, msg_to_bit_it_2_vnu_33_in_0, msg_to_bit_it_2_vnu_70_in_0, msg_to_bit_it_2_vnu_105_in_0, msg_to_bit_it_2_vnu_144_in_0, msg_to_bit_it_2_vnu_182_in_0);
cnu check_node_31_1(msg_to_check_it_1_cnu_31_in_0, msg_to_check_it_1_cnu_31_in_1, msg_to_check_it_1_cnu_31_in_2, msg_to_check_it_1_cnu_31_in_3, msg_to_check_it_1_cnu_31_in_4, msg_to_check_it_1_cnu_31_in_5, msg_to_bit_it_2_vnu_0_in_0, msg_to_bit_it_2_vnu_34_in_0, msg_to_bit_it_2_vnu_71_in_0, msg_to_bit_it_2_vnu_106_in_0, msg_to_bit_it_2_vnu_145_in_0, msg_to_bit_it_2_vnu_183_in_0);
cnu check_node_32_1(msg_to_check_it_1_cnu_32_in_0, msg_to_check_it_1_cnu_32_in_1, msg_to_check_it_1_cnu_32_in_2, msg_to_check_it_1_cnu_32_in_3, msg_to_check_it_1_cnu_32_in_4, msg_to_check_it_1_cnu_32_in_5, msg_to_bit_it_2_vnu_1_in_0, msg_to_bit_it_2_vnu_35_in_0, msg_to_bit_it_2_vnu_72_in_0, msg_to_bit_it_2_vnu_107_in_0, msg_to_bit_it_2_vnu_146_in_0, msg_to_bit_it_2_vnu_184_in_0);
cnu check_node_33_1(msg_to_check_it_1_cnu_33_in_0, msg_to_check_it_1_cnu_33_in_1, msg_to_check_it_1_cnu_33_in_2, msg_to_check_it_1_cnu_33_in_3, msg_to_check_it_1_cnu_33_in_4, msg_to_check_it_1_cnu_33_in_5, msg_to_bit_it_2_vnu_4_in_1, msg_to_bit_it_2_vnu_38_in_1, msg_to_bit_it_2_vnu_77_in_1, msg_to_bit_it_2_vnu_111_in_1, msg_to_bit_it_2_vnu_155_in_1, msg_to_bit_it_2_vnu_190_in_1);
cnu check_node_34_1(msg_to_check_it_1_cnu_34_in_0, msg_to_check_it_1_cnu_34_in_1, msg_to_check_it_1_cnu_34_in_2, msg_to_check_it_1_cnu_34_in_3, msg_to_check_it_1_cnu_34_in_4, msg_to_check_it_1_cnu_34_in_5, msg_to_bit_it_2_vnu_5_in_1, msg_to_bit_it_2_vnu_39_in_1, msg_to_bit_it_2_vnu_78_in_1, msg_to_bit_it_2_vnu_112_in_1, msg_to_bit_it_2_vnu_156_in_1, msg_to_bit_it_2_vnu_191_in_1);
cnu check_node_35_1(msg_to_check_it_1_cnu_35_in_0, msg_to_check_it_1_cnu_35_in_1, msg_to_check_it_1_cnu_35_in_2, msg_to_check_it_1_cnu_35_in_3, msg_to_check_it_1_cnu_35_in_4, msg_to_check_it_1_cnu_35_in_5, msg_to_bit_it_2_vnu_6_in_1, msg_to_bit_it_2_vnu_40_in_1, msg_to_bit_it_2_vnu_79_in_1, msg_to_bit_it_2_vnu_113_in_1, msg_to_bit_it_2_vnu_157_in_1, msg_to_bit_it_2_vnu_192_in_1);
cnu check_node_36_1(msg_to_check_it_1_cnu_36_in_0, msg_to_check_it_1_cnu_36_in_1, msg_to_check_it_1_cnu_36_in_2, msg_to_check_it_1_cnu_36_in_3, msg_to_check_it_1_cnu_36_in_4, msg_to_check_it_1_cnu_36_in_5, msg_to_bit_it_2_vnu_7_in_1, msg_to_bit_it_2_vnu_41_in_1, msg_to_bit_it_2_vnu_80_in_1, msg_to_bit_it_2_vnu_114_in_1, msg_to_bit_it_2_vnu_158_in_1, msg_to_bit_it_2_vnu_193_in_1);
cnu check_node_37_1(msg_to_check_it_1_cnu_37_in_0, msg_to_check_it_1_cnu_37_in_1, msg_to_check_it_1_cnu_37_in_2, msg_to_check_it_1_cnu_37_in_3, msg_to_check_it_1_cnu_37_in_4, msg_to_check_it_1_cnu_37_in_5, msg_to_bit_it_2_vnu_8_in_1, msg_to_bit_it_2_vnu_42_in_1, msg_to_bit_it_2_vnu_81_in_1, msg_to_bit_it_2_vnu_115_in_1, msg_to_bit_it_2_vnu_159_in_1, msg_to_bit_it_2_vnu_194_in_1);
cnu check_node_38_1(msg_to_check_it_1_cnu_38_in_0, msg_to_check_it_1_cnu_38_in_1, msg_to_check_it_1_cnu_38_in_2, msg_to_check_it_1_cnu_38_in_3, msg_to_check_it_1_cnu_38_in_4, msg_to_check_it_1_cnu_38_in_5, msg_to_bit_it_2_vnu_9_in_1, msg_to_bit_it_2_vnu_43_in_1, msg_to_bit_it_2_vnu_82_in_1, msg_to_bit_it_2_vnu_116_in_1, msg_to_bit_it_2_vnu_160_in_1, msg_to_bit_it_2_vnu_195_in_1);
cnu check_node_39_1(msg_to_check_it_1_cnu_39_in_0, msg_to_check_it_1_cnu_39_in_1, msg_to_check_it_1_cnu_39_in_2, msg_to_check_it_1_cnu_39_in_3, msg_to_check_it_1_cnu_39_in_4, msg_to_check_it_1_cnu_39_in_5, msg_to_bit_it_2_vnu_10_in_1, msg_to_bit_it_2_vnu_44_in_1, msg_to_bit_it_2_vnu_83_in_1, msg_to_bit_it_2_vnu_117_in_1, msg_to_bit_it_2_vnu_161_in_1, msg_to_bit_it_2_vnu_196_in_1);
cnu check_node_40_1(msg_to_check_it_1_cnu_40_in_0, msg_to_check_it_1_cnu_40_in_1, msg_to_check_it_1_cnu_40_in_2, msg_to_check_it_1_cnu_40_in_3, msg_to_check_it_1_cnu_40_in_4, msg_to_check_it_1_cnu_40_in_5, msg_to_bit_it_2_vnu_11_in_1, msg_to_bit_it_2_vnu_45_in_1, msg_to_bit_it_2_vnu_84_in_1, msg_to_bit_it_2_vnu_118_in_1, msg_to_bit_it_2_vnu_162_in_1, msg_to_bit_it_2_vnu_197_in_1);
cnu check_node_41_1(msg_to_check_it_1_cnu_41_in_0, msg_to_check_it_1_cnu_41_in_1, msg_to_check_it_1_cnu_41_in_2, msg_to_check_it_1_cnu_41_in_3, msg_to_check_it_1_cnu_41_in_4, msg_to_check_it_1_cnu_41_in_5, msg_to_bit_it_2_vnu_12_in_1, msg_to_bit_it_2_vnu_46_in_1, msg_to_bit_it_2_vnu_85_in_1, msg_to_bit_it_2_vnu_119_in_1, msg_to_bit_it_2_vnu_163_in_1, msg_to_bit_it_2_vnu_165_in_1);
cnu check_node_42_1(msg_to_check_it_1_cnu_42_in_0, msg_to_check_it_1_cnu_42_in_1, msg_to_check_it_1_cnu_42_in_2, msg_to_check_it_1_cnu_42_in_3, msg_to_check_it_1_cnu_42_in_4, msg_to_check_it_1_cnu_42_in_5, msg_to_bit_it_2_vnu_13_in_1, msg_to_bit_it_2_vnu_47_in_1, msg_to_bit_it_2_vnu_86_in_1, msg_to_bit_it_2_vnu_120_in_1, msg_to_bit_it_2_vnu_164_in_1, msg_to_bit_it_2_vnu_166_in_1);
cnu check_node_43_1(msg_to_check_it_1_cnu_43_in_0, msg_to_check_it_1_cnu_43_in_1, msg_to_check_it_1_cnu_43_in_2, msg_to_check_it_1_cnu_43_in_3, msg_to_check_it_1_cnu_43_in_4, msg_to_check_it_1_cnu_43_in_5, msg_to_bit_it_2_vnu_14_in_1, msg_to_bit_it_2_vnu_48_in_1, msg_to_bit_it_2_vnu_87_in_1, msg_to_bit_it_2_vnu_121_in_1, msg_to_bit_it_2_vnu_132_in_1, msg_to_bit_it_2_vnu_167_in_1);
cnu check_node_44_1(msg_to_check_it_1_cnu_44_in_0, msg_to_check_it_1_cnu_44_in_1, msg_to_check_it_1_cnu_44_in_2, msg_to_check_it_1_cnu_44_in_3, msg_to_check_it_1_cnu_44_in_4, msg_to_check_it_1_cnu_44_in_5, msg_to_bit_it_2_vnu_15_in_1, msg_to_bit_it_2_vnu_49_in_1, msg_to_bit_it_2_vnu_88_in_1, msg_to_bit_it_2_vnu_122_in_1, msg_to_bit_it_2_vnu_133_in_1, msg_to_bit_it_2_vnu_168_in_1);
cnu check_node_45_1(msg_to_check_it_1_cnu_45_in_0, msg_to_check_it_1_cnu_45_in_1, msg_to_check_it_1_cnu_45_in_2, msg_to_check_it_1_cnu_45_in_3, msg_to_check_it_1_cnu_45_in_4, msg_to_check_it_1_cnu_45_in_5, msg_to_bit_it_2_vnu_16_in_1, msg_to_bit_it_2_vnu_50_in_1, msg_to_bit_it_2_vnu_89_in_1, msg_to_bit_it_2_vnu_123_in_1, msg_to_bit_it_2_vnu_134_in_1, msg_to_bit_it_2_vnu_169_in_1);
cnu check_node_46_1(msg_to_check_it_1_cnu_46_in_0, msg_to_check_it_1_cnu_46_in_1, msg_to_check_it_1_cnu_46_in_2, msg_to_check_it_1_cnu_46_in_3, msg_to_check_it_1_cnu_46_in_4, msg_to_check_it_1_cnu_46_in_5, msg_to_bit_it_2_vnu_17_in_1, msg_to_bit_it_2_vnu_51_in_1, msg_to_bit_it_2_vnu_90_in_1, msg_to_bit_it_2_vnu_124_in_1, msg_to_bit_it_2_vnu_135_in_1, msg_to_bit_it_2_vnu_170_in_1);
cnu check_node_47_1(msg_to_check_it_1_cnu_47_in_0, msg_to_check_it_1_cnu_47_in_1, msg_to_check_it_1_cnu_47_in_2, msg_to_check_it_1_cnu_47_in_3, msg_to_check_it_1_cnu_47_in_4, msg_to_check_it_1_cnu_47_in_5, msg_to_bit_it_2_vnu_18_in_1, msg_to_bit_it_2_vnu_52_in_1, msg_to_bit_it_2_vnu_91_in_1, msg_to_bit_it_2_vnu_125_in_1, msg_to_bit_it_2_vnu_136_in_1, msg_to_bit_it_2_vnu_171_in_1);
cnu check_node_48_1(msg_to_check_it_1_cnu_48_in_0, msg_to_check_it_1_cnu_48_in_1, msg_to_check_it_1_cnu_48_in_2, msg_to_check_it_1_cnu_48_in_3, msg_to_check_it_1_cnu_48_in_4, msg_to_check_it_1_cnu_48_in_5, msg_to_bit_it_2_vnu_19_in_1, msg_to_bit_it_2_vnu_53_in_1, msg_to_bit_it_2_vnu_92_in_1, msg_to_bit_it_2_vnu_126_in_1, msg_to_bit_it_2_vnu_137_in_1, msg_to_bit_it_2_vnu_172_in_1);
cnu check_node_49_1(msg_to_check_it_1_cnu_49_in_0, msg_to_check_it_1_cnu_49_in_1, msg_to_check_it_1_cnu_49_in_2, msg_to_check_it_1_cnu_49_in_3, msg_to_check_it_1_cnu_49_in_4, msg_to_check_it_1_cnu_49_in_5, msg_to_bit_it_2_vnu_20_in_1, msg_to_bit_it_2_vnu_54_in_1, msg_to_bit_it_2_vnu_93_in_1, msg_to_bit_it_2_vnu_127_in_1, msg_to_bit_it_2_vnu_138_in_1, msg_to_bit_it_2_vnu_173_in_1);
cnu check_node_50_1(msg_to_check_it_1_cnu_50_in_0, msg_to_check_it_1_cnu_50_in_1, msg_to_check_it_1_cnu_50_in_2, msg_to_check_it_1_cnu_50_in_3, msg_to_check_it_1_cnu_50_in_4, msg_to_check_it_1_cnu_50_in_5, msg_to_bit_it_2_vnu_21_in_1, msg_to_bit_it_2_vnu_55_in_1, msg_to_bit_it_2_vnu_94_in_1, msg_to_bit_it_2_vnu_128_in_1, msg_to_bit_it_2_vnu_139_in_1, msg_to_bit_it_2_vnu_174_in_1);
cnu check_node_51_1(msg_to_check_it_1_cnu_51_in_0, msg_to_check_it_1_cnu_51_in_1, msg_to_check_it_1_cnu_51_in_2, msg_to_check_it_1_cnu_51_in_3, msg_to_check_it_1_cnu_51_in_4, msg_to_check_it_1_cnu_51_in_5, msg_to_bit_it_2_vnu_22_in_1, msg_to_bit_it_2_vnu_56_in_1, msg_to_bit_it_2_vnu_95_in_1, msg_to_bit_it_2_vnu_129_in_1, msg_to_bit_it_2_vnu_140_in_1, msg_to_bit_it_2_vnu_175_in_1);
cnu check_node_52_1(msg_to_check_it_1_cnu_52_in_0, msg_to_check_it_1_cnu_52_in_1, msg_to_check_it_1_cnu_52_in_2, msg_to_check_it_1_cnu_52_in_3, msg_to_check_it_1_cnu_52_in_4, msg_to_check_it_1_cnu_52_in_5, msg_to_bit_it_2_vnu_23_in_1, msg_to_bit_it_2_vnu_57_in_1, msg_to_bit_it_2_vnu_96_in_1, msg_to_bit_it_2_vnu_130_in_1, msg_to_bit_it_2_vnu_141_in_1, msg_to_bit_it_2_vnu_176_in_1);
cnu check_node_53_1(msg_to_check_it_1_cnu_53_in_0, msg_to_check_it_1_cnu_53_in_1, msg_to_check_it_1_cnu_53_in_2, msg_to_check_it_1_cnu_53_in_3, msg_to_check_it_1_cnu_53_in_4, msg_to_check_it_1_cnu_53_in_5, msg_to_bit_it_2_vnu_24_in_1, msg_to_bit_it_2_vnu_58_in_1, msg_to_bit_it_2_vnu_97_in_1, msg_to_bit_it_2_vnu_131_in_1, msg_to_bit_it_2_vnu_142_in_1, msg_to_bit_it_2_vnu_177_in_1);
cnu check_node_54_1(msg_to_check_it_1_cnu_54_in_0, msg_to_check_it_1_cnu_54_in_1, msg_to_check_it_1_cnu_54_in_2, msg_to_check_it_1_cnu_54_in_3, msg_to_check_it_1_cnu_54_in_4, msg_to_check_it_1_cnu_54_in_5, msg_to_bit_it_2_vnu_25_in_1, msg_to_bit_it_2_vnu_59_in_1, msg_to_bit_it_2_vnu_98_in_1, msg_to_bit_it_2_vnu_99_in_1, msg_to_bit_it_2_vnu_143_in_1, msg_to_bit_it_2_vnu_178_in_1);
cnu check_node_55_1(msg_to_check_it_1_cnu_55_in_0, msg_to_check_it_1_cnu_55_in_1, msg_to_check_it_1_cnu_55_in_2, msg_to_check_it_1_cnu_55_in_3, msg_to_check_it_1_cnu_55_in_4, msg_to_check_it_1_cnu_55_in_5, msg_to_bit_it_2_vnu_26_in_1, msg_to_bit_it_2_vnu_60_in_1, msg_to_bit_it_2_vnu_66_in_1, msg_to_bit_it_2_vnu_100_in_1, msg_to_bit_it_2_vnu_144_in_1, msg_to_bit_it_2_vnu_179_in_1);
cnu check_node_56_1(msg_to_check_it_1_cnu_56_in_0, msg_to_check_it_1_cnu_56_in_1, msg_to_check_it_1_cnu_56_in_2, msg_to_check_it_1_cnu_56_in_3, msg_to_check_it_1_cnu_56_in_4, msg_to_check_it_1_cnu_56_in_5, msg_to_bit_it_2_vnu_27_in_1, msg_to_bit_it_2_vnu_61_in_1, msg_to_bit_it_2_vnu_67_in_1, msg_to_bit_it_2_vnu_101_in_1, msg_to_bit_it_2_vnu_145_in_1, msg_to_bit_it_2_vnu_180_in_1);
cnu check_node_57_1(msg_to_check_it_1_cnu_57_in_0, msg_to_check_it_1_cnu_57_in_1, msg_to_check_it_1_cnu_57_in_2, msg_to_check_it_1_cnu_57_in_3, msg_to_check_it_1_cnu_57_in_4, msg_to_check_it_1_cnu_57_in_5, msg_to_bit_it_2_vnu_28_in_1, msg_to_bit_it_2_vnu_62_in_1, msg_to_bit_it_2_vnu_68_in_1, msg_to_bit_it_2_vnu_102_in_1, msg_to_bit_it_2_vnu_146_in_1, msg_to_bit_it_2_vnu_181_in_1);
cnu check_node_58_1(msg_to_check_it_1_cnu_58_in_0, msg_to_check_it_1_cnu_58_in_1, msg_to_check_it_1_cnu_58_in_2, msg_to_check_it_1_cnu_58_in_3, msg_to_check_it_1_cnu_58_in_4, msg_to_check_it_1_cnu_58_in_5, msg_to_bit_it_2_vnu_29_in_1, msg_to_bit_it_2_vnu_63_in_1, msg_to_bit_it_2_vnu_69_in_1, msg_to_bit_it_2_vnu_103_in_1, msg_to_bit_it_2_vnu_147_in_1, msg_to_bit_it_2_vnu_182_in_1);
cnu check_node_59_1(msg_to_check_it_1_cnu_59_in_0, msg_to_check_it_1_cnu_59_in_1, msg_to_check_it_1_cnu_59_in_2, msg_to_check_it_1_cnu_59_in_3, msg_to_check_it_1_cnu_59_in_4, msg_to_check_it_1_cnu_59_in_5, msg_to_bit_it_2_vnu_30_in_1, msg_to_bit_it_2_vnu_64_in_1, msg_to_bit_it_2_vnu_70_in_1, msg_to_bit_it_2_vnu_104_in_1, msg_to_bit_it_2_vnu_148_in_1, msg_to_bit_it_2_vnu_183_in_1);
cnu check_node_60_1(msg_to_check_it_1_cnu_60_in_0, msg_to_check_it_1_cnu_60_in_1, msg_to_check_it_1_cnu_60_in_2, msg_to_check_it_1_cnu_60_in_3, msg_to_check_it_1_cnu_60_in_4, msg_to_check_it_1_cnu_60_in_5, msg_to_bit_it_2_vnu_31_in_1, msg_to_bit_it_2_vnu_65_in_1, msg_to_bit_it_2_vnu_71_in_1, msg_to_bit_it_2_vnu_105_in_1, msg_to_bit_it_2_vnu_149_in_1, msg_to_bit_it_2_vnu_184_in_1);
cnu check_node_61_1(msg_to_check_it_1_cnu_61_in_0, msg_to_check_it_1_cnu_61_in_1, msg_to_check_it_1_cnu_61_in_2, msg_to_check_it_1_cnu_61_in_3, msg_to_check_it_1_cnu_61_in_4, msg_to_check_it_1_cnu_61_in_5, msg_to_bit_it_2_vnu_32_in_1, msg_to_bit_it_2_vnu_33_in_1, msg_to_bit_it_2_vnu_72_in_1, msg_to_bit_it_2_vnu_106_in_1, msg_to_bit_it_2_vnu_150_in_1, msg_to_bit_it_2_vnu_185_in_1);
cnu check_node_62_1(msg_to_check_it_1_cnu_62_in_0, msg_to_check_it_1_cnu_62_in_1, msg_to_check_it_1_cnu_62_in_2, msg_to_check_it_1_cnu_62_in_3, msg_to_check_it_1_cnu_62_in_4, msg_to_check_it_1_cnu_62_in_5, msg_to_bit_it_2_vnu_0_in_1, msg_to_bit_it_2_vnu_34_in_1, msg_to_bit_it_2_vnu_73_in_1, msg_to_bit_it_2_vnu_107_in_1, msg_to_bit_it_2_vnu_151_in_1, msg_to_bit_it_2_vnu_186_in_1);
cnu check_node_63_1(msg_to_check_it_1_cnu_63_in_0, msg_to_check_it_1_cnu_63_in_1, msg_to_check_it_1_cnu_63_in_2, msg_to_check_it_1_cnu_63_in_3, msg_to_check_it_1_cnu_63_in_4, msg_to_check_it_1_cnu_63_in_5, msg_to_bit_it_2_vnu_1_in_1, msg_to_bit_it_2_vnu_35_in_1, msg_to_bit_it_2_vnu_74_in_1, msg_to_bit_it_2_vnu_108_in_1, msg_to_bit_it_2_vnu_152_in_1, msg_to_bit_it_2_vnu_187_in_1);
cnu check_node_64_1(msg_to_check_it_1_cnu_64_in_0, msg_to_check_it_1_cnu_64_in_1, msg_to_check_it_1_cnu_64_in_2, msg_to_check_it_1_cnu_64_in_3, msg_to_check_it_1_cnu_64_in_4, msg_to_check_it_1_cnu_64_in_5, msg_to_bit_it_2_vnu_2_in_1, msg_to_bit_it_2_vnu_36_in_1, msg_to_bit_it_2_vnu_75_in_1, msg_to_bit_it_2_vnu_109_in_1, msg_to_bit_it_2_vnu_153_in_1, msg_to_bit_it_2_vnu_188_in_1);
cnu check_node_65_1(msg_to_check_it_1_cnu_65_in_0, msg_to_check_it_1_cnu_65_in_1, msg_to_check_it_1_cnu_65_in_2, msg_to_check_it_1_cnu_65_in_3, msg_to_check_it_1_cnu_65_in_4, msg_to_check_it_1_cnu_65_in_5, msg_to_bit_it_2_vnu_3_in_1, msg_to_bit_it_2_vnu_37_in_1, msg_to_bit_it_2_vnu_76_in_1, msg_to_bit_it_2_vnu_110_in_1, msg_to_bit_it_2_vnu_154_in_1, msg_to_bit_it_2_vnu_189_in_1);
cnu check_node_66_1(msg_to_check_it_1_cnu_66_in_0, msg_to_check_it_1_cnu_66_in_1, msg_to_check_it_1_cnu_66_in_2, msg_to_check_it_1_cnu_66_in_3, msg_to_check_it_1_cnu_66_in_4, msg_to_check_it_1_cnu_66_in_5, msg_to_bit_it_2_vnu_6_in_2, msg_to_bit_it_2_vnu_41_in_2, msg_to_bit_it_2_vnu_80_in_2, msg_to_bit_it_2_vnu_118_in_2, msg_to_bit_it_2_vnu_159_in_2, msg_to_bit_it_2_vnu_195_in_2);
cnu check_node_67_1(msg_to_check_it_1_cnu_67_in_0, msg_to_check_it_1_cnu_67_in_1, msg_to_check_it_1_cnu_67_in_2, msg_to_check_it_1_cnu_67_in_3, msg_to_check_it_1_cnu_67_in_4, msg_to_check_it_1_cnu_67_in_5, msg_to_bit_it_2_vnu_7_in_2, msg_to_bit_it_2_vnu_42_in_2, msg_to_bit_it_2_vnu_81_in_2, msg_to_bit_it_2_vnu_119_in_2, msg_to_bit_it_2_vnu_160_in_2, msg_to_bit_it_2_vnu_196_in_2);
cnu check_node_68_1(msg_to_check_it_1_cnu_68_in_0, msg_to_check_it_1_cnu_68_in_1, msg_to_check_it_1_cnu_68_in_2, msg_to_check_it_1_cnu_68_in_3, msg_to_check_it_1_cnu_68_in_4, msg_to_check_it_1_cnu_68_in_5, msg_to_bit_it_2_vnu_8_in_2, msg_to_bit_it_2_vnu_43_in_2, msg_to_bit_it_2_vnu_82_in_2, msg_to_bit_it_2_vnu_120_in_2, msg_to_bit_it_2_vnu_161_in_2, msg_to_bit_it_2_vnu_197_in_2);
cnu check_node_69_1(msg_to_check_it_1_cnu_69_in_0, msg_to_check_it_1_cnu_69_in_1, msg_to_check_it_1_cnu_69_in_2, msg_to_check_it_1_cnu_69_in_3, msg_to_check_it_1_cnu_69_in_4, msg_to_check_it_1_cnu_69_in_5, msg_to_bit_it_2_vnu_9_in_2, msg_to_bit_it_2_vnu_44_in_2, msg_to_bit_it_2_vnu_83_in_2, msg_to_bit_it_2_vnu_121_in_2, msg_to_bit_it_2_vnu_162_in_2, msg_to_bit_it_2_vnu_165_in_2);
cnu check_node_70_1(msg_to_check_it_1_cnu_70_in_0, msg_to_check_it_1_cnu_70_in_1, msg_to_check_it_1_cnu_70_in_2, msg_to_check_it_1_cnu_70_in_3, msg_to_check_it_1_cnu_70_in_4, msg_to_check_it_1_cnu_70_in_5, msg_to_bit_it_2_vnu_10_in_2, msg_to_bit_it_2_vnu_45_in_2, msg_to_bit_it_2_vnu_84_in_2, msg_to_bit_it_2_vnu_122_in_2, msg_to_bit_it_2_vnu_163_in_2, msg_to_bit_it_2_vnu_166_in_2);
cnu check_node_71_1(msg_to_check_it_1_cnu_71_in_0, msg_to_check_it_1_cnu_71_in_1, msg_to_check_it_1_cnu_71_in_2, msg_to_check_it_1_cnu_71_in_3, msg_to_check_it_1_cnu_71_in_4, msg_to_check_it_1_cnu_71_in_5, msg_to_bit_it_2_vnu_11_in_2, msg_to_bit_it_2_vnu_46_in_2, msg_to_bit_it_2_vnu_85_in_2, msg_to_bit_it_2_vnu_123_in_2, msg_to_bit_it_2_vnu_164_in_2, msg_to_bit_it_2_vnu_167_in_2);
cnu check_node_72_1(msg_to_check_it_1_cnu_72_in_0, msg_to_check_it_1_cnu_72_in_1, msg_to_check_it_1_cnu_72_in_2, msg_to_check_it_1_cnu_72_in_3, msg_to_check_it_1_cnu_72_in_4, msg_to_check_it_1_cnu_72_in_5, msg_to_bit_it_2_vnu_12_in_2, msg_to_bit_it_2_vnu_47_in_2, msg_to_bit_it_2_vnu_86_in_2, msg_to_bit_it_2_vnu_124_in_2, msg_to_bit_it_2_vnu_132_in_2, msg_to_bit_it_2_vnu_168_in_2);
cnu check_node_73_1(msg_to_check_it_1_cnu_73_in_0, msg_to_check_it_1_cnu_73_in_1, msg_to_check_it_1_cnu_73_in_2, msg_to_check_it_1_cnu_73_in_3, msg_to_check_it_1_cnu_73_in_4, msg_to_check_it_1_cnu_73_in_5, msg_to_bit_it_2_vnu_13_in_2, msg_to_bit_it_2_vnu_48_in_2, msg_to_bit_it_2_vnu_87_in_2, msg_to_bit_it_2_vnu_125_in_2, msg_to_bit_it_2_vnu_133_in_2, msg_to_bit_it_2_vnu_169_in_2);
cnu check_node_74_1(msg_to_check_it_1_cnu_74_in_0, msg_to_check_it_1_cnu_74_in_1, msg_to_check_it_1_cnu_74_in_2, msg_to_check_it_1_cnu_74_in_3, msg_to_check_it_1_cnu_74_in_4, msg_to_check_it_1_cnu_74_in_5, msg_to_bit_it_2_vnu_14_in_2, msg_to_bit_it_2_vnu_49_in_2, msg_to_bit_it_2_vnu_88_in_2, msg_to_bit_it_2_vnu_126_in_2, msg_to_bit_it_2_vnu_134_in_2, msg_to_bit_it_2_vnu_170_in_2);
cnu check_node_75_1(msg_to_check_it_1_cnu_75_in_0, msg_to_check_it_1_cnu_75_in_1, msg_to_check_it_1_cnu_75_in_2, msg_to_check_it_1_cnu_75_in_3, msg_to_check_it_1_cnu_75_in_4, msg_to_check_it_1_cnu_75_in_5, msg_to_bit_it_2_vnu_15_in_2, msg_to_bit_it_2_vnu_50_in_2, msg_to_bit_it_2_vnu_89_in_2, msg_to_bit_it_2_vnu_127_in_2, msg_to_bit_it_2_vnu_135_in_2, msg_to_bit_it_2_vnu_171_in_2);
cnu check_node_76_1(msg_to_check_it_1_cnu_76_in_0, msg_to_check_it_1_cnu_76_in_1, msg_to_check_it_1_cnu_76_in_2, msg_to_check_it_1_cnu_76_in_3, msg_to_check_it_1_cnu_76_in_4, msg_to_check_it_1_cnu_76_in_5, msg_to_bit_it_2_vnu_16_in_2, msg_to_bit_it_2_vnu_51_in_2, msg_to_bit_it_2_vnu_90_in_2, msg_to_bit_it_2_vnu_128_in_2, msg_to_bit_it_2_vnu_136_in_2, msg_to_bit_it_2_vnu_172_in_2);
cnu check_node_77_1(msg_to_check_it_1_cnu_77_in_0, msg_to_check_it_1_cnu_77_in_1, msg_to_check_it_1_cnu_77_in_2, msg_to_check_it_1_cnu_77_in_3, msg_to_check_it_1_cnu_77_in_4, msg_to_check_it_1_cnu_77_in_5, msg_to_bit_it_2_vnu_17_in_2, msg_to_bit_it_2_vnu_52_in_2, msg_to_bit_it_2_vnu_91_in_2, msg_to_bit_it_2_vnu_129_in_2, msg_to_bit_it_2_vnu_137_in_2, msg_to_bit_it_2_vnu_173_in_2);
cnu check_node_78_1(msg_to_check_it_1_cnu_78_in_0, msg_to_check_it_1_cnu_78_in_1, msg_to_check_it_1_cnu_78_in_2, msg_to_check_it_1_cnu_78_in_3, msg_to_check_it_1_cnu_78_in_4, msg_to_check_it_1_cnu_78_in_5, msg_to_bit_it_2_vnu_18_in_2, msg_to_bit_it_2_vnu_53_in_2, msg_to_bit_it_2_vnu_92_in_2, msg_to_bit_it_2_vnu_130_in_2, msg_to_bit_it_2_vnu_138_in_2, msg_to_bit_it_2_vnu_174_in_2);
cnu check_node_79_1(msg_to_check_it_1_cnu_79_in_0, msg_to_check_it_1_cnu_79_in_1, msg_to_check_it_1_cnu_79_in_2, msg_to_check_it_1_cnu_79_in_3, msg_to_check_it_1_cnu_79_in_4, msg_to_check_it_1_cnu_79_in_5, msg_to_bit_it_2_vnu_19_in_2, msg_to_bit_it_2_vnu_54_in_2, msg_to_bit_it_2_vnu_93_in_2, msg_to_bit_it_2_vnu_131_in_2, msg_to_bit_it_2_vnu_139_in_2, msg_to_bit_it_2_vnu_175_in_2);
cnu check_node_80_1(msg_to_check_it_1_cnu_80_in_0, msg_to_check_it_1_cnu_80_in_1, msg_to_check_it_1_cnu_80_in_2, msg_to_check_it_1_cnu_80_in_3, msg_to_check_it_1_cnu_80_in_4, msg_to_check_it_1_cnu_80_in_5, msg_to_bit_it_2_vnu_20_in_2, msg_to_bit_it_2_vnu_55_in_2, msg_to_bit_it_2_vnu_94_in_2, msg_to_bit_it_2_vnu_99_in_2, msg_to_bit_it_2_vnu_140_in_2, msg_to_bit_it_2_vnu_176_in_2);
cnu check_node_81_1(msg_to_check_it_1_cnu_81_in_0, msg_to_check_it_1_cnu_81_in_1, msg_to_check_it_1_cnu_81_in_2, msg_to_check_it_1_cnu_81_in_3, msg_to_check_it_1_cnu_81_in_4, msg_to_check_it_1_cnu_81_in_5, msg_to_bit_it_2_vnu_21_in_2, msg_to_bit_it_2_vnu_56_in_2, msg_to_bit_it_2_vnu_95_in_2, msg_to_bit_it_2_vnu_100_in_2, msg_to_bit_it_2_vnu_141_in_2, msg_to_bit_it_2_vnu_177_in_2);
cnu check_node_82_1(msg_to_check_it_1_cnu_82_in_0, msg_to_check_it_1_cnu_82_in_1, msg_to_check_it_1_cnu_82_in_2, msg_to_check_it_1_cnu_82_in_3, msg_to_check_it_1_cnu_82_in_4, msg_to_check_it_1_cnu_82_in_5, msg_to_bit_it_2_vnu_22_in_2, msg_to_bit_it_2_vnu_57_in_2, msg_to_bit_it_2_vnu_96_in_2, msg_to_bit_it_2_vnu_101_in_2, msg_to_bit_it_2_vnu_142_in_2, msg_to_bit_it_2_vnu_178_in_2);
cnu check_node_83_1(msg_to_check_it_1_cnu_83_in_0, msg_to_check_it_1_cnu_83_in_1, msg_to_check_it_1_cnu_83_in_2, msg_to_check_it_1_cnu_83_in_3, msg_to_check_it_1_cnu_83_in_4, msg_to_check_it_1_cnu_83_in_5, msg_to_bit_it_2_vnu_23_in_2, msg_to_bit_it_2_vnu_58_in_2, msg_to_bit_it_2_vnu_97_in_2, msg_to_bit_it_2_vnu_102_in_2, msg_to_bit_it_2_vnu_143_in_2, msg_to_bit_it_2_vnu_179_in_2);
cnu check_node_84_1(msg_to_check_it_1_cnu_84_in_0, msg_to_check_it_1_cnu_84_in_1, msg_to_check_it_1_cnu_84_in_2, msg_to_check_it_1_cnu_84_in_3, msg_to_check_it_1_cnu_84_in_4, msg_to_check_it_1_cnu_84_in_5, msg_to_bit_it_2_vnu_24_in_2, msg_to_bit_it_2_vnu_59_in_2, msg_to_bit_it_2_vnu_98_in_2, msg_to_bit_it_2_vnu_103_in_2, msg_to_bit_it_2_vnu_144_in_2, msg_to_bit_it_2_vnu_180_in_2);
cnu check_node_85_1(msg_to_check_it_1_cnu_85_in_0, msg_to_check_it_1_cnu_85_in_1, msg_to_check_it_1_cnu_85_in_2, msg_to_check_it_1_cnu_85_in_3, msg_to_check_it_1_cnu_85_in_4, msg_to_check_it_1_cnu_85_in_5, msg_to_bit_it_2_vnu_25_in_2, msg_to_bit_it_2_vnu_60_in_2, msg_to_bit_it_2_vnu_66_in_2, msg_to_bit_it_2_vnu_104_in_2, msg_to_bit_it_2_vnu_145_in_2, msg_to_bit_it_2_vnu_181_in_2);
cnu check_node_86_1(msg_to_check_it_1_cnu_86_in_0, msg_to_check_it_1_cnu_86_in_1, msg_to_check_it_1_cnu_86_in_2, msg_to_check_it_1_cnu_86_in_3, msg_to_check_it_1_cnu_86_in_4, msg_to_check_it_1_cnu_86_in_5, msg_to_bit_it_2_vnu_26_in_2, msg_to_bit_it_2_vnu_61_in_2, msg_to_bit_it_2_vnu_67_in_2, msg_to_bit_it_2_vnu_105_in_2, msg_to_bit_it_2_vnu_146_in_2, msg_to_bit_it_2_vnu_182_in_2);
cnu check_node_87_1(msg_to_check_it_1_cnu_87_in_0, msg_to_check_it_1_cnu_87_in_1, msg_to_check_it_1_cnu_87_in_2, msg_to_check_it_1_cnu_87_in_3, msg_to_check_it_1_cnu_87_in_4, msg_to_check_it_1_cnu_87_in_5, msg_to_bit_it_2_vnu_27_in_2, msg_to_bit_it_2_vnu_62_in_2, msg_to_bit_it_2_vnu_68_in_2, msg_to_bit_it_2_vnu_106_in_2, msg_to_bit_it_2_vnu_147_in_2, msg_to_bit_it_2_vnu_183_in_2);
cnu check_node_88_1(msg_to_check_it_1_cnu_88_in_0, msg_to_check_it_1_cnu_88_in_1, msg_to_check_it_1_cnu_88_in_2, msg_to_check_it_1_cnu_88_in_3, msg_to_check_it_1_cnu_88_in_4, msg_to_check_it_1_cnu_88_in_5, msg_to_bit_it_2_vnu_28_in_2, msg_to_bit_it_2_vnu_63_in_2, msg_to_bit_it_2_vnu_69_in_2, msg_to_bit_it_2_vnu_107_in_2, msg_to_bit_it_2_vnu_148_in_2, msg_to_bit_it_2_vnu_184_in_2);
cnu check_node_89_1(msg_to_check_it_1_cnu_89_in_0, msg_to_check_it_1_cnu_89_in_1, msg_to_check_it_1_cnu_89_in_2, msg_to_check_it_1_cnu_89_in_3, msg_to_check_it_1_cnu_89_in_4, msg_to_check_it_1_cnu_89_in_5, msg_to_bit_it_2_vnu_29_in_2, msg_to_bit_it_2_vnu_64_in_2, msg_to_bit_it_2_vnu_70_in_2, msg_to_bit_it_2_vnu_108_in_2, msg_to_bit_it_2_vnu_149_in_2, msg_to_bit_it_2_vnu_185_in_2);
cnu check_node_90_1(msg_to_check_it_1_cnu_90_in_0, msg_to_check_it_1_cnu_90_in_1, msg_to_check_it_1_cnu_90_in_2, msg_to_check_it_1_cnu_90_in_3, msg_to_check_it_1_cnu_90_in_4, msg_to_check_it_1_cnu_90_in_5, msg_to_bit_it_2_vnu_30_in_2, msg_to_bit_it_2_vnu_65_in_2, msg_to_bit_it_2_vnu_71_in_2, msg_to_bit_it_2_vnu_109_in_2, msg_to_bit_it_2_vnu_150_in_2, msg_to_bit_it_2_vnu_186_in_2);
cnu check_node_91_1(msg_to_check_it_1_cnu_91_in_0, msg_to_check_it_1_cnu_91_in_1, msg_to_check_it_1_cnu_91_in_2, msg_to_check_it_1_cnu_91_in_3, msg_to_check_it_1_cnu_91_in_4, msg_to_check_it_1_cnu_91_in_5, msg_to_bit_it_2_vnu_31_in_2, msg_to_bit_it_2_vnu_33_in_2, msg_to_bit_it_2_vnu_72_in_2, msg_to_bit_it_2_vnu_110_in_2, msg_to_bit_it_2_vnu_151_in_2, msg_to_bit_it_2_vnu_187_in_2);
cnu check_node_92_1(msg_to_check_it_1_cnu_92_in_0, msg_to_check_it_1_cnu_92_in_1, msg_to_check_it_1_cnu_92_in_2, msg_to_check_it_1_cnu_92_in_3, msg_to_check_it_1_cnu_92_in_4, msg_to_check_it_1_cnu_92_in_5, msg_to_bit_it_2_vnu_32_in_2, msg_to_bit_it_2_vnu_34_in_2, msg_to_bit_it_2_vnu_73_in_2, msg_to_bit_it_2_vnu_111_in_2, msg_to_bit_it_2_vnu_152_in_2, msg_to_bit_it_2_vnu_188_in_2);
cnu check_node_93_1(msg_to_check_it_1_cnu_93_in_0, msg_to_check_it_1_cnu_93_in_1, msg_to_check_it_1_cnu_93_in_2, msg_to_check_it_1_cnu_93_in_3, msg_to_check_it_1_cnu_93_in_4, msg_to_check_it_1_cnu_93_in_5, msg_to_bit_it_2_vnu_0_in_2, msg_to_bit_it_2_vnu_35_in_2, msg_to_bit_it_2_vnu_74_in_2, msg_to_bit_it_2_vnu_112_in_2, msg_to_bit_it_2_vnu_153_in_2, msg_to_bit_it_2_vnu_189_in_2);
cnu check_node_94_1(msg_to_check_it_1_cnu_94_in_0, msg_to_check_it_1_cnu_94_in_1, msg_to_check_it_1_cnu_94_in_2, msg_to_check_it_1_cnu_94_in_3, msg_to_check_it_1_cnu_94_in_4, msg_to_check_it_1_cnu_94_in_5, msg_to_bit_it_2_vnu_1_in_2, msg_to_bit_it_2_vnu_36_in_2, msg_to_bit_it_2_vnu_75_in_2, msg_to_bit_it_2_vnu_113_in_2, msg_to_bit_it_2_vnu_154_in_2, msg_to_bit_it_2_vnu_190_in_2);
cnu check_node_95_1(msg_to_check_it_1_cnu_95_in_0, msg_to_check_it_1_cnu_95_in_1, msg_to_check_it_1_cnu_95_in_2, msg_to_check_it_1_cnu_95_in_3, msg_to_check_it_1_cnu_95_in_4, msg_to_check_it_1_cnu_95_in_5, msg_to_bit_it_2_vnu_2_in_2, msg_to_bit_it_2_vnu_37_in_2, msg_to_bit_it_2_vnu_76_in_2, msg_to_bit_it_2_vnu_114_in_2, msg_to_bit_it_2_vnu_155_in_2, msg_to_bit_it_2_vnu_191_in_2);
cnu check_node_96_1(msg_to_check_it_1_cnu_96_in_0, msg_to_check_it_1_cnu_96_in_1, msg_to_check_it_1_cnu_96_in_2, msg_to_check_it_1_cnu_96_in_3, msg_to_check_it_1_cnu_96_in_4, msg_to_check_it_1_cnu_96_in_5, msg_to_bit_it_2_vnu_3_in_2, msg_to_bit_it_2_vnu_38_in_2, msg_to_bit_it_2_vnu_77_in_2, msg_to_bit_it_2_vnu_115_in_2, msg_to_bit_it_2_vnu_156_in_2, msg_to_bit_it_2_vnu_192_in_2);
cnu check_node_97_1(msg_to_check_it_1_cnu_97_in_0, msg_to_check_it_1_cnu_97_in_1, msg_to_check_it_1_cnu_97_in_2, msg_to_check_it_1_cnu_97_in_3, msg_to_check_it_1_cnu_97_in_4, msg_to_check_it_1_cnu_97_in_5, msg_to_bit_it_2_vnu_4_in_2, msg_to_bit_it_2_vnu_39_in_2, msg_to_bit_it_2_vnu_78_in_2, msg_to_bit_it_2_vnu_116_in_2, msg_to_bit_it_2_vnu_157_in_2, msg_to_bit_it_2_vnu_193_in_2);
cnu check_node_98_1(msg_to_check_it_1_cnu_98_in_0, msg_to_check_it_1_cnu_98_in_1, msg_to_check_it_1_cnu_98_in_2, msg_to_check_it_1_cnu_98_in_3, msg_to_check_it_1_cnu_98_in_4, msg_to_check_it_1_cnu_98_in_5, msg_to_bit_it_2_vnu_5_in_2, msg_to_bit_it_2_vnu_40_in_2, msg_to_bit_it_2_vnu_79_in_2, msg_to_bit_it_2_vnu_117_in_2, msg_to_bit_it_2_vnu_158_in_2, msg_to_bit_it_2_vnu_194_in_2);


vnu_h hard_dec0(data_0, msg_to_bit_it_2_vnu_0_in_0, msg_to_bit_it_2_vnu_0_in_1, msg_to_bit_it_2_vnu_0_in_2, data_out[0]);
vnu_h hard_dec1(data_1, msg_to_bit_it_2_vnu_1_in_0, msg_to_bit_it_2_vnu_1_in_1, msg_to_bit_it_2_vnu_1_in_2, data_out[1]);
vnu_h hard_dec2(data_2, msg_to_bit_it_2_vnu_2_in_0, msg_to_bit_it_2_vnu_2_in_1, msg_to_bit_it_2_vnu_2_in_2, data_out[2]);
vnu_h hard_dec3(data_3, msg_to_bit_it_2_vnu_3_in_0, msg_to_bit_it_2_vnu_3_in_1, msg_to_bit_it_2_vnu_3_in_2, data_out[3]);
vnu_h hard_dec4(data_4, msg_to_bit_it_2_vnu_4_in_0, msg_to_bit_it_2_vnu_4_in_1, msg_to_bit_it_2_vnu_4_in_2, data_out[4]);
vnu_h hard_dec5(data_5, msg_to_bit_it_2_vnu_5_in_0, msg_to_bit_it_2_vnu_5_in_1, msg_to_bit_it_2_vnu_5_in_2, data_out[5]);
vnu_h hard_dec6(data_6, msg_to_bit_it_2_vnu_6_in_0, msg_to_bit_it_2_vnu_6_in_1, msg_to_bit_it_2_vnu_6_in_2, data_out[6]);
vnu_h hard_dec7(data_7, msg_to_bit_it_2_vnu_7_in_0, msg_to_bit_it_2_vnu_7_in_1, msg_to_bit_it_2_vnu_7_in_2, data_out[7]);
vnu_h hard_dec8(data_8, msg_to_bit_it_2_vnu_8_in_0, msg_to_bit_it_2_vnu_8_in_1, msg_to_bit_it_2_vnu_8_in_2, data_out[8]);
vnu_h hard_dec9(data_9, msg_to_bit_it_2_vnu_9_in_0, msg_to_bit_it_2_vnu_9_in_1, msg_to_bit_it_2_vnu_9_in_2, data_out[9]);
vnu_h hard_dec10(data_10, msg_to_bit_it_2_vnu_10_in_0, msg_to_bit_it_2_vnu_10_in_1, msg_to_bit_it_2_vnu_10_in_2, data_out[10]);
vnu_h hard_dec11(data_11, msg_to_bit_it_2_vnu_11_in_0, msg_to_bit_it_2_vnu_11_in_1, msg_to_bit_it_2_vnu_11_in_2, data_out[11]);
vnu_h hard_dec12(data_12, msg_to_bit_it_2_vnu_12_in_0, msg_to_bit_it_2_vnu_12_in_1, msg_to_bit_it_2_vnu_12_in_2, data_out[12]);
vnu_h hard_dec13(data_13, msg_to_bit_it_2_vnu_13_in_0, msg_to_bit_it_2_vnu_13_in_1, msg_to_bit_it_2_vnu_13_in_2, data_out[13]);
vnu_h hard_dec14(data_14, msg_to_bit_it_2_vnu_14_in_0, msg_to_bit_it_2_vnu_14_in_1, msg_to_bit_it_2_vnu_14_in_2, data_out[14]);
vnu_h hard_dec15(data_15, msg_to_bit_it_2_vnu_15_in_0, msg_to_bit_it_2_vnu_15_in_1, msg_to_bit_it_2_vnu_15_in_2, data_out[15]);
vnu_h hard_dec16(data_16, msg_to_bit_it_2_vnu_16_in_0, msg_to_bit_it_2_vnu_16_in_1, msg_to_bit_it_2_vnu_16_in_2, data_out[16]);
vnu_h hard_dec17(data_17, msg_to_bit_it_2_vnu_17_in_0, msg_to_bit_it_2_vnu_17_in_1, msg_to_bit_it_2_vnu_17_in_2, data_out[17]);
vnu_h hard_dec18(data_18, msg_to_bit_it_2_vnu_18_in_0, msg_to_bit_it_2_vnu_18_in_1, msg_to_bit_it_2_vnu_18_in_2, data_out[18]);
vnu_h hard_dec19(data_19, msg_to_bit_it_2_vnu_19_in_0, msg_to_bit_it_2_vnu_19_in_1, msg_to_bit_it_2_vnu_19_in_2, data_out[19]);
vnu_h hard_dec20(data_20, msg_to_bit_it_2_vnu_20_in_0, msg_to_bit_it_2_vnu_20_in_1, msg_to_bit_it_2_vnu_20_in_2, data_out[20]);
vnu_h hard_dec21(data_21, msg_to_bit_it_2_vnu_21_in_0, msg_to_bit_it_2_vnu_21_in_1, msg_to_bit_it_2_vnu_21_in_2, data_out[21]);
vnu_h hard_dec22(data_22, msg_to_bit_it_2_vnu_22_in_0, msg_to_bit_it_2_vnu_22_in_1, msg_to_bit_it_2_vnu_22_in_2, data_out[22]);
vnu_h hard_dec23(data_23, msg_to_bit_it_2_vnu_23_in_0, msg_to_bit_it_2_vnu_23_in_1, msg_to_bit_it_2_vnu_23_in_2, data_out[23]);
vnu_h hard_dec24(data_24, msg_to_bit_it_2_vnu_24_in_0, msg_to_bit_it_2_vnu_24_in_1, msg_to_bit_it_2_vnu_24_in_2, data_out[24]);
vnu_h hard_dec25(data_25, msg_to_bit_it_2_vnu_25_in_0, msg_to_bit_it_2_vnu_25_in_1, msg_to_bit_it_2_vnu_25_in_2, data_out[25]);
vnu_h hard_dec26(data_26, msg_to_bit_it_2_vnu_26_in_0, msg_to_bit_it_2_vnu_26_in_1, msg_to_bit_it_2_vnu_26_in_2, data_out[26]);
vnu_h hard_dec27(data_27, msg_to_bit_it_2_vnu_27_in_0, msg_to_bit_it_2_vnu_27_in_1, msg_to_bit_it_2_vnu_27_in_2, data_out[27]);
vnu_h hard_dec28(data_28, msg_to_bit_it_2_vnu_28_in_0, msg_to_bit_it_2_vnu_28_in_1, msg_to_bit_it_2_vnu_28_in_2, data_out[28]);
vnu_h hard_dec29(data_29, msg_to_bit_it_2_vnu_29_in_0, msg_to_bit_it_2_vnu_29_in_1, msg_to_bit_it_2_vnu_29_in_2, data_out[29]);
vnu_h hard_dec30(data_30, msg_to_bit_it_2_vnu_30_in_0, msg_to_bit_it_2_vnu_30_in_1, msg_to_bit_it_2_vnu_30_in_2, data_out[30]);
vnu_h hard_dec31(data_31, msg_to_bit_it_2_vnu_31_in_0, msg_to_bit_it_2_vnu_31_in_1, msg_to_bit_it_2_vnu_31_in_2, data_out[31]);
vnu_h hard_dec32(data_32, msg_to_bit_it_2_vnu_32_in_0, msg_to_bit_it_2_vnu_32_in_1, msg_to_bit_it_2_vnu_32_in_2, data_out[32]);
vnu_h hard_dec33(data_33, msg_to_bit_it_2_vnu_33_in_0, msg_to_bit_it_2_vnu_33_in_1, msg_to_bit_it_2_vnu_33_in_2, data_out[33]);
vnu_h hard_dec34(data_34, msg_to_bit_it_2_vnu_34_in_0, msg_to_bit_it_2_vnu_34_in_1, msg_to_bit_it_2_vnu_34_in_2, data_out[34]);
vnu_h hard_dec35(data_35, msg_to_bit_it_2_vnu_35_in_0, msg_to_bit_it_2_vnu_35_in_1, msg_to_bit_it_2_vnu_35_in_2, data_out[35]);
vnu_h hard_dec36(data_36, msg_to_bit_it_2_vnu_36_in_0, msg_to_bit_it_2_vnu_36_in_1, msg_to_bit_it_2_vnu_36_in_2, data_out[36]);
vnu_h hard_dec37(data_37, msg_to_bit_it_2_vnu_37_in_0, msg_to_bit_it_2_vnu_37_in_1, msg_to_bit_it_2_vnu_37_in_2, data_out[37]);
vnu_h hard_dec38(data_38, msg_to_bit_it_2_vnu_38_in_0, msg_to_bit_it_2_vnu_38_in_1, msg_to_bit_it_2_vnu_38_in_2, data_out[38]);
vnu_h hard_dec39(data_39, msg_to_bit_it_2_vnu_39_in_0, msg_to_bit_it_2_vnu_39_in_1, msg_to_bit_it_2_vnu_39_in_2, data_out[39]);
vnu_h hard_dec40(data_40, msg_to_bit_it_2_vnu_40_in_0, msg_to_bit_it_2_vnu_40_in_1, msg_to_bit_it_2_vnu_40_in_2, data_out[40]);
vnu_h hard_dec41(data_41, msg_to_bit_it_2_vnu_41_in_0, msg_to_bit_it_2_vnu_41_in_1, msg_to_bit_it_2_vnu_41_in_2, data_out[41]);
vnu_h hard_dec42(data_42, msg_to_bit_it_2_vnu_42_in_0, msg_to_bit_it_2_vnu_42_in_1, msg_to_bit_it_2_vnu_42_in_2, data_out[42]);
vnu_h hard_dec43(data_43, msg_to_bit_it_2_vnu_43_in_0, msg_to_bit_it_2_vnu_43_in_1, msg_to_bit_it_2_vnu_43_in_2, data_out[43]);
vnu_h hard_dec44(data_44, msg_to_bit_it_2_vnu_44_in_0, msg_to_bit_it_2_vnu_44_in_1, msg_to_bit_it_2_vnu_44_in_2, data_out[44]);
vnu_h hard_dec45(data_45, msg_to_bit_it_2_vnu_45_in_0, msg_to_bit_it_2_vnu_45_in_1, msg_to_bit_it_2_vnu_45_in_2, data_out[45]);
vnu_h hard_dec46(data_46, msg_to_bit_it_2_vnu_46_in_0, msg_to_bit_it_2_vnu_46_in_1, msg_to_bit_it_2_vnu_46_in_2, data_out[46]);
vnu_h hard_dec47(data_47, msg_to_bit_it_2_vnu_47_in_0, msg_to_bit_it_2_vnu_47_in_1, msg_to_bit_it_2_vnu_47_in_2, data_out[47]);
vnu_h hard_dec48(data_48, msg_to_bit_it_2_vnu_48_in_0, msg_to_bit_it_2_vnu_48_in_1, msg_to_bit_it_2_vnu_48_in_2, data_out[48]);
vnu_h hard_dec49(data_49, msg_to_bit_it_2_vnu_49_in_0, msg_to_bit_it_2_vnu_49_in_1, msg_to_bit_it_2_vnu_49_in_2, data_out[49]);
vnu_h hard_dec50(data_50, msg_to_bit_it_2_vnu_50_in_0, msg_to_bit_it_2_vnu_50_in_1, msg_to_bit_it_2_vnu_50_in_2, data_out[50]);
vnu_h hard_dec51(data_51, msg_to_bit_it_2_vnu_51_in_0, msg_to_bit_it_2_vnu_51_in_1, msg_to_bit_it_2_vnu_51_in_2, data_out[51]);
vnu_h hard_dec52(data_52, msg_to_bit_it_2_vnu_52_in_0, msg_to_bit_it_2_vnu_52_in_1, msg_to_bit_it_2_vnu_52_in_2, data_out[52]);
vnu_h hard_dec53(data_53, msg_to_bit_it_2_vnu_53_in_0, msg_to_bit_it_2_vnu_53_in_1, msg_to_bit_it_2_vnu_53_in_2, data_out[53]);
vnu_h hard_dec54(data_54, msg_to_bit_it_2_vnu_54_in_0, msg_to_bit_it_2_vnu_54_in_1, msg_to_bit_it_2_vnu_54_in_2, data_out[54]);
vnu_h hard_dec55(data_55, msg_to_bit_it_2_vnu_55_in_0, msg_to_bit_it_2_vnu_55_in_1, msg_to_bit_it_2_vnu_55_in_2, data_out[55]);
vnu_h hard_dec56(data_56, msg_to_bit_it_2_vnu_56_in_0, msg_to_bit_it_2_vnu_56_in_1, msg_to_bit_it_2_vnu_56_in_2, data_out[56]);
vnu_h hard_dec57(data_57, msg_to_bit_it_2_vnu_57_in_0, msg_to_bit_it_2_vnu_57_in_1, msg_to_bit_it_2_vnu_57_in_2, data_out[57]);
vnu_h hard_dec58(data_58, msg_to_bit_it_2_vnu_58_in_0, msg_to_bit_it_2_vnu_58_in_1, msg_to_bit_it_2_vnu_58_in_2, data_out[58]);
vnu_h hard_dec59(data_59, msg_to_bit_it_2_vnu_59_in_0, msg_to_bit_it_2_vnu_59_in_1, msg_to_bit_it_2_vnu_59_in_2, data_out[59]);
vnu_h hard_dec60(data_60, msg_to_bit_it_2_vnu_60_in_0, msg_to_bit_it_2_vnu_60_in_1, msg_to_bit_it_2_vnu_60_in_2, data_out[60]);
vnu_h hard_dec61(data_61, msg_to_bit_it_2_vnu_61_in_0, msg_to_bit_it_2_vnu_61_in_1, msg_to_bit_it_2_vnu_61_in_2, data_out[61]);
vnu_h hard_dec62(data_62, msg_to_bit_it_2_vnu_62_in_0, msg_to_bit_it_2_vnu_62_in_1, msg_to_bit_it_2_vnu_62_in_2, data_out[62]);
vnu_h hard_dec63(data_63, msg_to_bit_it_2_vnu_63_in_0, msg_to_bit_it_2_vnu_63_in_1, msg_to_bit_it_2_vnu_63_in_2, data_out[63]);
vnu_h hard_dec64(data_64, msg_to_bit_it_2_vnu_64_in_0, msg_to_bit_it_2_vnu_64_in_1, msg_to_bit_it_2_vnu_64_in_2, data_out[64]);
vnu_h hard_dec65(data_65, msg_to_bit_it_2_vnu_65_in_0, msg_to_bit_it_2_vnu_65_in_1, msg_to_bit_it_2_vnu_65_in_2, data_out[65]);
vnu_h hard_dec66(data_66, msg_to_bit_it_2_vnu_66_in_0, msg_to_bit_it_2_vnu_66_in_1, msg_to_bit_it_2_vnu_66_in_2, data_out[66]);
vnu_h hard_dec67(data_67, msg_to_bit_it_2_vnu_67_in_0, msg_to_bit_it_2_vnu_67_in_1, msg_to_bit_it_2_vnu_67_in_2, data_out[67]);
vnu_h hard_dec68(data_68, msg_to_bit_it_2_vnu_68_in_0, msg_to_bit_it_2_vnu_68_in_1, msg_to_bit_it_2_vnu_68_in_2, data_out[68]);
vnu_h hard_dec69(data_69, msg_to_bit_it_2_vnu_69_in_0, msg_to_bit_it_2_vnu_69_in_1, msg_to_bit_it_2_vnu_69_in_2, data_out[69]);
vnu_h hard_dec70(data_70, msg_to_bit_it_2_vnu_70_in_0, msg_to_bit_it_2_vnu_70_in_1, msg_to_bit_it_2_vnu_70_in_2, data_out[70]);
vnu_h hard_dec71(data_71, msg_to_bit_it_2_vnu_71_in_0, msg_to_bit_it_2_vnu_71_in_1, msg_to_bit_it_2_vnu_71_in_2, data_out[71]);
vnu_h hard_dec72(data_72, msg_to_bit_it_2_vnu_72_in_0, msg_to_bit_it_2_vnu_72_in_1, msg_to_bit_it_2_vnu_72_in_2, data_out[72]);
vnu_h hard_dec73(data_73, msg_to_bit_it_2_vnu_73_in_0, msg_to_bit_it_2_vnu_73_in_1, msg_to_bit_it_2_vnu_73_in_2, data_out[73]);
vnu_h hard_dec74(data_74, msg_to_bit_it_2_vnu_74_in_0, msg_to_bit_it_2_vnu_74_in_1, msg_to_bit_it_2_vnu_74_in_2, data_out[74]);
vnu_h hard_dec75(data_75, msg_to_bit_it_2_vnu_75_in_0, msg_to_bit_it_2_vnu_75_in_1, msg_to_bit_it_2_vnu_75_in_2, data_out[75]);
vnu_h hard_dec76(data_76, msg_to_bit_it_2_vnu_76_in_0, msg_to_bit_it_2_vnu_76_in_1, msg_to_bit_it_2_vnu_76_in_2, data_out[76]);
vnu_h hard_dec77(data_77, msg_to_bit_it_2_vnu_77_in_0, msg_to_bit_it_2_vnu_77_in_1, msg_to_bit_it_2_vnu_77_in_2, data_out[77]);
vnu_h hard_dec78(data_78, msg_to_bit_it_2_vnu_78_in_0, msg_to_bit_it_2_vnu_78_in_1, msg_to_bit_it_2_vnu_78_in_2, data_out[78]);
vnu_h hard_dec79(data_79, msg_to_bit_it_2_vnu_79_in_0, msg_to_bit_it_2_vnu_79_in_1, msg_to_bit_it_2_vnu_79_in_2, data_out[79]);
vnu_h hard_dec80(data_80, msg_to_bit_it_2_vnu_80_in_0, msg_to_bit_it_2_vnu_80_in_1, msg_to_bit_it_2_vnu_80_in_2, data_out[80]);
vnu_h hard_dec81(data_81, msg_to_bit_it_2_vnu_81_in_0, msg_to_bit_it_2_vnu_81_in_1, msg_to_bit_it_2_vnu_81_in_2, data_out[81]);
vnu_h hard_dec82(data_82, msg_to_bit_it_2_vnu_82_in_0, msg_to_bit_it_2_vnu_82_in_1, msg_to_bit_it_2_vnu_82_in_2, data_out[82]);
vnu_h hard_dec83(data_83, msg_to_bit_it_2_vnu_83_in_0, msg_to_bit_it_2_vnu_83_in_1, msg_to_bit_it_2_vnu_83_in_2, data_out[83]);
vnu_h hard_dec84(data_84, msg_to_bit_it_2_vnu_84_in_0, msg_to_bit_it_2_vnu_84_in_1, msg_to_bit_it_2_vnu_84_in_2, data_out[84]);
vnu_h hard_dec85(data_85, msg_to_bit_it_2_vnu_85_in_0, msg_to_bit_it_2_vnu_85_in_1, msg_to_bit_it_2_vnu_85_in_2, data_out[85]);
vnu_h hard_dec86(data_86, msg_to_bit_it_2_vnu_86_in_0, msg_to_bit_it_2_vnu_86_in_1, msg_to_bit_it_2_vnu_86_in_2, data_out[86]);
vnu_h hard_dec87(data_87, msg_to_bit_it_2_vnu_87_in_0, msg_to_bit_it_2_vnu_87_in_1, msg_to_bit_it_2_vnu_87_in_2, data_out[87]);
vnu_h hard_dec88(data_88, msg_to_bit_it_2_vnu_88_in_0, msg_to_bit_it_2_vnu_88_in_1, msg_to_bit_it_2_vnu_88_in_2, data_out[88]);
vnu_h hard_dec89(data_89, msg_to_bit_it_2_vnu_89_in_0, msg_to_bit_it_2_vnu_89_in_1, msg_to_bit_it_2_vnu_89_in_2, data_out[89]);
vnu_h hard_dec90(data_90, msg_to_bit_it_2_vnu_90_in_0, msg_to_bit_it_2_vnu_90_in_1, msg_to_bit_it_2_vnu_90_in_2, data_out[90]);
vnu_h hard_dec91(data_91, msg_to_bit_it_2_vnu_91_in_0, msg_to_bit_it_2_vnu_91_in_1, msg_to_bit_it_2_vnu_91_in_2, data_out[91]);
vnu_h hard_dec92(data_92, msg_to_bit_it_2_vnu_92_in_0, msg_to_bit_it_2_vnu_92_in_1, msg_to_bit_it_2_vnu_92_in_2, data_out[92]);
vnu_h hard_dec93(data_93, msg_to_bit_it_2_vnu_93_in_0, msg_to_bit_it_2_vnu_93_in_1, msg_to_bit_it_2_vnu_93_in_2, data_out[93]);
vnu_h hard_dec94(data_94, msg_to_bit_it_2_vnu_94_in_0, msg_to_bit_it_2_vnu_94_in_1, msg_to_bit_it_2_vnu_94_in_2, data_out[94]);
vnu_h hard_dec95(data_95, msg_to_bit_it_2_vnu_95_in_0, msg_to_bit_it_2_vnu_95_in_1, msg_to_bit_it_2_vnu_95_in_2, data_out[95]);
vnu_h hard_dec96(data_96, msg_to_bit_it_2_vnu_96_in_0, msg_to_bit_it_2_vnu_96_in_1, msg_to_bit_it_2_vnu_96_in_2, data_out[96]);
vnu_h hard_dec97(data_97, msg_to_bit_it_2_vnu_97_in_0, msg_to_bit_it_2_vnu_97_in_1, msg_to_bit_it_2_vnu_97_in_2, data_out[97]);
vnu_h hard_dec98(data_98, msg_to_bit_it_2_vnu_98_in_0, msg_to_bit_it_2_vnu_98_in_1, msg_to_bit_it_2_vnu_98_in_2, data_out[98]);
vnu_h hard_dec99(data_99, msg_to_bit_it_2_vnu_99_in_0, msg_to_bit_it_2_vnu_99_in_1, msg_to_bit_it_2_vnu_99_in_2, data_out[99]);
vnu_h hard_dec100(data_100, msg_to_bit_it_2_vnu_100_in_0, msg_to_bit_it_2_vnu_100_in_1, msg_to_bit_it_2_vnu_100_in_2, data_out[100]);
vnu_h hard_dec101(data_101, msg_to_bit_it_2_vnu_101_in_0, msg_to_bit_it_2_vnu_101_in_1, msg_to_bit_it_2_vnu_101_in_2, data_out[101]);
vnu_h hard_dec102(data_102, msg_to_bit_it_2_vnu_102_in_0, msg_to_bit_it_2_vnu_102_in_1, msg_to_bit_it_2_vnu_102_in_2, data_out[102]);
vnu_h hard_dec103(data_103, msg_to_bit_it_2_vnu_103_in_0, msg_to_bit_it_2_vnu_103_in_1, msg_to_bit_it_2_vnu_103_in_2, data_out[103]);
vnu_h hard_dec104(data_104, msg_to_bit_it_2_vnu_104_in_0, msg_to_bit_it_2_vnu_104_in_1, msg_to_bit_it_2_vnu_104_in_2, data_out[104]);
vnu_h hard_dec105(data_105, msg_to_bit_it_2_vnu_105_in_0, msg_to_bit_it_2_vnu_105_in_1, msg_to_bit_it_2_vnu_105_in_2, data_out[105]);
vnu_h hard_dec106(data_106, msg_to_bit_it_2_vnu_106_in_0, msg_to_bit_it_2_vnu_106_in_1, msg_to_bit_it_2_vnu_106_in_2, data_out[106]);
vnu_h hard_dec107(data_107, msg_to_bit_it_2_vnu_107_in_0, msg_to_bit_it_2_vnu_107_in_1, msg_to_bit_it_2_vnu_107_in_2, data_out[107]);
vnu_h hard_dec108(data_108, msg_to_bit_it_2_vnu_108_in_0, msg_to_bit_it_2_vnu_108_in_1, msg_to_bit_it_2_vnu_108_in_2, data_out[108]);
vnu_h hard_dec109(data_109, msg_to_bit_it_2_vnu_109_in_0, msg_to_bit_it_2_vnu_109_in_1, msg_to_bit_it_2_vnu_109_in_2, data_out[109]);
vnu_h hard_dec110(data_110, msg_to_bit_it_2_vnu_110_in_0, msg_to_bit_it_2_vnu_110_in_1, msg_to_bit_it_2_vnu_110_in_2, data_out[110]);
vnu_h hard_dec111(data_111, msg_to_bit_it_2_vnu_111_in_0, msg_to_bit_it_2_vnu_111_in_1, msg_to_bit_it_2_vnu_111_in_2, data_out[111]);
vnu_h hard_dec112(data_112, msg_to_bit_it_2_vnu_112_in_0, msg_to_bit_it_2_vnu_112_in_1, msg_to_bit_it_2_vnu_112_in_2, data_out[112]);
vnu_h hard_dec113(data_113, msg_to_bit_it_2_vnu_113_in_0, msg_to_bit_it_2_vnu_113_in_1, msg_to_bit_it_2_vnu_113_in_2, data_out[113]);
vnu_h hard_dec114(data_114, msg_to_bit_it_2_vnu_114_in_0, msg_to_bit_it_2_vnu_114_in_1, msg_to_bit_it_2_vnu_114_in_2, data_out[114]);
vnu_h hard_dec115(data_115, msg_to_bit_it_2_vnu_115_in_0, msg_to_bit_it_2_vnu_115_in_1, msg_to_bit_it_2_vnu_115_in_2, data_out[115]);
vnu_h hard_dec116(data_116, msg_to_bit_it_2_vnu_116_in_0, msg_to_bit_it_2_vnu_116_in_1, msg_to_bit_it_2_vnu_116_in_2, data_out[116]);
vnu_h hard_dec117(data_117, msg_to_bit_it_2_vnu_117_in_0, msg_to_bit_it_2_vnu_117_in_1, msg_to_bit_it_2_vnu_117_in_2, data_out[117]);
vnu_h hard_dec118(data_118, msg_to_bit_it_2_vnu_118_in_0, msg_to_bit_it_2_vnu_118_in_1, msg_to_bit_it_2_vnu_118_in_2, data_out[118]);
vnu_h hard_dec119(data_119, msg_to_bit_it_2_vnu_119_in_0, msg_to_bit_it_2_vnu_119_in_1, msg_to_bit_it_2_vnu_119_in_2, data_out[119]);
vnu_h hard_dec120(data_120, msg_to_bit_it_2_vnu_120_in_0, msg_to_bit_it_2_vnu_120_in_1, msg_to_bit_it_2_vnu_120_in_2, data_out[120]);
vnu_h hard_dec121(data_121, msg_to_bit_it_2_vnu_121_in_0, msg_to_bit_it_2_vnu_121_in_1, msg_to_bit_it_2_vnu_121_in_2, data_out[121]);
vnu_h hard_dec122(data_122, msg_to_bit_it_2_vnu_122_in_0, msg_to_bit_it_2_vnu_122_in_1, msg_to_bit_it_2_vnu_122_in_2, data_out[122]);
vnu_h hard_dec123(data_123, msg_to_bit_it_2_vnu_123_in_0, msg_to_bit_it_2_vnu_123_in_1, msg_to_bit_it_2_vnu_123_in_2, data_out[123]);
vnu_h hard_dec124(data_124, msg_to_bit_it_2_vnu_124_in_0, msg_to_bit_it_2_vnu_124_in_1, msg_to_bit_it_2_vnu_124_in_2, data_out[124]);
vnu_h hard_dec125(data_125, msg_to_bit_it_2_vnu_125_in_0, msg_to_bit_it_2_vnu_125_in_1, msg_to_bit_it_2_vnu_125_in_2, data_out[125]);
vnu_h hard_dec126(data_126, msg_to_bit_it_2_vnu_126_in_0, msg_to_bit_it_2_vnu_126_in_1, msg_to_bit_it_2_vnu_126_in_2, data_out[126]);
vnu_h hard_dec127(data_127, msg_to_bit_it_2_vnu_127_in_0, msg_to_bit_it_2_vnu_127_in_1, msg_to_bit_it_2_vnu_127_in_2, data_out[127]);
vnu_h hard_dec128(data_128, msg_to_bit_it_2_vnu_128_in_0, msg_to_bit_it_2_vnu_128_in_1, msg_to_bit_it_2_vnu_128_in_2, data_out[128]);
vnu_h hard_dec129(data_129, msg_to_bit_it_2_vnu_129_in_0, msg_to_bit_it_2_vnu_129_in_1, msg_to_bit_it_2_vnu_129_in_2, data_out[129]);
vnu_h hard_dec130(data_130, msg_to_bit_it_2_vnu_130_in_0, msg_to_bit_it_2_vnu_130_in_1, msg_to_bit_it_2_vnu_130_in_2, data_out[130]);
vnu_h hard_dec131(data_131, msg_to_bit_it_2_vnu_131_in_0, msg_to_bit_it_2_vnu_131_in_1, msg_to_bit_it_2_vnu_131_in_2, data_out[131]);
vnu_h hard_dec132(data_132, msg_to_bit_it_2_vnu_132_in_0, msg_to_bit_it_2_vnu_132_in_1, msg_to_bit_it_2_vnu_132_in_2, data_out[132]);
vnu_h hard_dec133(data_133, msg_to_bit_it_2_vnu_133_in_0, msg_to_bit_it_2_vnu_133_in_1, msg_to_bit_it_2_vnu_133_in_2, data_out[133]);
vnu_h hard_dec134(data_134, msg_to_bit_it_2_vnu_134_in_0, msg_to_bit_it_2_vnu_134_in_1, msg_to_bit_it_2_vnu_134_in_2, data_out[134]);
vnu_h hard_dec135(data_135, msg_to_bit_it_2_vnu_135_in_0, msg_to_bit_it_2_vnu_135_in_1, msg_to_bit_it_2_vnu_135_in_2, data_out[135]);
vnu_h hard_dec136(data_136, msg_to_bit_it_2_vnu_136_in_0, msg_to_bit_it_2_vnu_136_in_1, msg_to_bit_it_2_vnu_136_in_2, data_out[136]);
vnu_h hard_dec137(data_137, msg_to_bit_it_2_vnu_137_in_0, msg_to_bit_it_2_vnu_137_in_1, msg_to_bit_it_2_vnu_137_in_2, data_out[137]);
vnu_h hard_dec138(data_138, msg_to_bit_it_2_vnu_138_in_0, msg_to_bit_it_2_vnu_138_in_1, msg_to_bit_it_2_vnu_138_in_2, data_out[138]);
vnu_h hard_dec139(data_139, msg_to_bit_it_2_vnu_139_in_0, msg_to_bit_it_2_vnu_139_in_1, msg_to_bit_it_2_vnu_139_in_2, data_out[139]);
vnu_h hard_dec140(data_140, msg_to_bit_it_2_vnu_140_in_0, msg_to_bit_it_2_vnu_140_in_1, msg_to_bit_it_2_vnu_140_in_2, data_out[140]);
vnu_h hard_dec141(data_141, msg_to_bit_it_2_vnu_141_in_0, msg_to_bit_it_2_vnu_141_in_1, msg_to_bit_it_2_vnu_141_in_2, data_out[141]);
vnu_h hard_dec142(data_142, msg_to_bit_it_2_vnu_142_in_0, msg_to_bit_it_2_vnu_142_in_1, msg_to_bit_it_2_vnu_142_in_2, data_out[142]);
vnu_h hard_dec143(data_143, msg_to_bit_it_2_vnu_143_in_0, msg_to_bit_it_2_vnu_143_in_1, msg_to_bit_it_2_vnu_143_in_2, data_out[143]);
vnu_h hard_dec144(data_144, msg_to_bit_it_2_vnu_144_in_0, msg_to_bit_it_2_vnu_144_in_1, msg_to_bit_it_2_vnu_144_in_2, data_out[144]);
vnu_h hard_dec145(data_145, msg_to_bit_it_2_vnu_145_in_0, msg_to_bit_it_2_vnu_145_in_1, msg_to_bit_it_2_vnu_145_in_2, data_out[145]);
vnu_h hard_dec146(data_146, msg_to_bit_it_2_vnu_146_in_0, msg_to_bit_it_2_vnu_146_in_1, msg_to_bit_it_2_vnu_146_in_2, data_out[146]);
vnu_h hard_dec147(data_147, msg_to_bit_it_2_vnu_147_in_0, msg_to_bit_it_2_vnu_147_in_1, msg_to_bit_it_2_vnu_147_in_2, data_out[147]);
vnu_h hard_dec148(data_148, msg_to_bit_it_2_vnu_148_in_0, msg_to_bit_it_2_vnu_148_in_1, msg_to_bit_it_2_vnu_148_in_2, data_out[148]);
vnu_h hard_dec149(data_149, msg_to_bit_it_2_vnu_149_in_0, msg_to_bit_it_2_vnu_149_in_1, msg_to_bit_it_2_vnu_149_in_2, data_out[149]);
vnu_h hard_dec150(data_150, msg_to_bit_it_2_vnu_150_in_0, msg_to_bit_it_2_vnu_150_in_1, msg_to_bit_it_2_vnu_150_in_2, data_out[150]);
vnu_h hard_dec151(data_151, msg_to_bit_it_2_vnu_151_in_0, msg_to_bit_it_2_vnu_151_in_1, msg_to_bit_it_2_vnu_151_in_2, data_out[151]);
vnu_h hard_dec152(data_152, msg_to_bit_it_2_vnu_152_in_0, msg_to_bit_it_2_vnu_152_in_1, msg_to_bit_it_2_vnu_152_in_2, data_out[152]);
vnu_h hard_dec153(data_153, msg_to_bit_it_2_vnu_153_in_0, msg_to_bit_it_2_vnu_153_in_1, msg_to_bit_it_2_vnu_153_in_2, data_out[153]);
vnu_h hard_dec154(data_154, msg_to_bit_it_2_vnu_154_in_0, msg_to_bit_it_2_vnu_154_in_1, msg_to_bit_it_2_vnu_154_in_2, data_out[154]);
vnu_h hard_dec155(data_155, msg_to_bit_it_2_vnu_155_in_0, msg_to_bit_it_2_vnu_155_in_1, msg_to_bit_it_2_vnu_155_in_2, data_out[155]);
vnu_h hard_dec156(data_156, msg_to_bit_it_2_vnu_156_in_0, msg_to_bit_it_2_vnu_156_in_1, msg_to_bit_it_2_vnu_156_in_2, data_out[156]);
vnu_h hard_dec157(data_157, msg_to_bit_it_2_vnu_157_in_0, msg_to_bit_it_2_vnu_157_in_1, msg_to_bit_it_2_vnu_157_in_2, data_out[157]);
vnu_h hard_dec158(data_158, msg_to_bit_it_2_vnu_158_in_0, msg_to_bit_it_2_vnu_158_in_1, msg_to_bit_it_2_vnu_158_in_2, data_out[158]);
vnu_h hard_dec159(data_159, msg_to_bit_it_2_vnu_159_in_0, msg_to_bit_it_2_vnu_159_in_1, msg_to_bit_it_2_vnu_159_in_2, data_out[159]);
vnu_h hard_dec160(data_160, msg_to_bit_it_2_vnu_160_in_0, msg_to_bit_it_2_vnu_160_in_1, msg_to_bit_it_2_vnu_160_in_2, data_out[160]);
vnu_h hard_dec161(data_161, msg_to_bit_it_2_vnu_161_in_0, msg_to_bit_it_2_vnu_161_in_1, msg_to_bit_it_2_vnu_161_in_2, data_out[161]);
vnu_h hard_dec162(data_162, msg_to_bit_it_2_vnu_162_in_0, msg_to_bit_it_2_vnu_162_in_1, msg_to_bit_it_2_vnu_162_in_2, data_out[162]);
vnu_h hard_dec163(data_163, msg_to_bit_it_2_vnu_163_in_0, msg_to_bit_it_2_vnu_163_in_1, msg_to_bit_it_2_vnu_163_in_2, data_out[163]);
vnu_h hard_dec164(data_164, msg_to_bit_it_2_vnu_164_in_0, msg_to_bit_it_2_vnu_164_in_1, msg_to_bit_it_2_vnu_164_in_2, data_out[164]);
vnu_h hard_dec165(data_165, msg_to_bit_it_2_vnu_165_in_0, msg_to_bit_it_2_vnu_165_in_1, msg_to_bit_it_2_vnu_165_in_2, data_out[165]);
vnu_h hard_dec166(data_166, msg_to_bit_it_2_vnu_166_in_0, msg_to_bit_it_2_vnu_166_in_1, msg_to_bit_it_2_vnu_166_in_2, data_out[166]);
vnu_h hard_dec167(data_167, msg_to_bit_it_2_vnu_167_in_0, msg_to_bit_it_2_vnu_167_in_1, msg_to_bit_it_2_vnu_167_in_2, data_out[167]);
vnu_h hard_dec168(data_168, msg_to_bit_it_2_vnu_168_in_0, msg_to_bit_it_2_vnu_168_in_1, msg_to_bit_it_2_vnu_168_in_2, data_out[168]);
vnu_h hard_dec169(data_169, msg_to_bit_it_2_vnu_169_in_0, msg_to_bit_it_2_vnu_169_in_1, msg_to_bit_it_2_vnu_169_in_2, data_out[169]);
vnu_h hard_dec170(data_170, msg_to_bit_it_2_vnu_170_in_0, msg_to_bit_it_2_vnu_170_in_1, msg_to_bit_it_2_vnu_170_in_2, data_out[170]);
vnu_h hard_dec171(data_171, msg_to_bit_it_2_vnu_171_in_0, msg_to_bit_it_2_vnu_171_in_1, msg_to_bit_it_2_vnu_171_in_2, data_out[171]);
vnu_h hard_dec172(data_172, msg_to_bit_it_2_vnu_172_in_0, msg_to_bit_it_2_vnu_172_in_1, msg_to_bit_it_2_vnu_172_in_2, data_out[172]);
vnu_h hard_dec173(data_173, msg_to_bit_it_2_vnu_173_in_0, msg_to_bit_it_2_vnu_173_in_1, msg_to_bit_it_2_vnu_173_in_2, data_out[173]);
vnu_h hard_dec174(data_174, msg_to_bit_it_2_vnu_174_in_0, msg_to_bit_it_2_vnu_174_in_1, msg_to_bit_it_2_vnu_174_in_2, data_out[174]);
vnu_h hard_dec175(data_175, msg_to_bit_it_2_vnu_175_in_0, msg_to_bit_it_2_vnu_175_in_1, msg_to_bit_it_2_vnu_175_in_2, data_out[175]);
vnu_h hard_dec176(data_176, msg_to_bit_it_2_vnu_176_in_0, msg_to_bit_it_2_vnu_176_in_1, msg_to_bit_it_2_vnu_176_in_2, data_out[176]);
vnu_h hard_dec177(data_177, msg_to_bit_it_2_vnu_177_in_0, msg_to_bit_it_2_vnu_177_in_1, msg_to_bit_it_2_vnu_177_in_2, data_out[177]);
vnu_h hard_dec178(data_178, msg_to_bit_it_2_vnu_178_in_0, msg_to_bit_it_2_vnu_178_in_1, msg_to_bit_it_2_vnu_178_in_2, data_out[178]);
vnu_h hard_dec179(data_179, msg_to_bit_it_2_vnu_179_in_0, msg_to_bit_it_2_vnu_179_in_1, msg_to_bit_it_2_vnu_179_in_2, data_out[179]);
vnu_h hard_dec180(data_180, msg_to_bit_it_2_vnu_180_in_0, msg_to_bit_it_2_vnu_180_in_1, msg_to_bit_it_2_vnu_180_in_2, data_out[180]);
vnu_h hard_dec181(data_181, msg_to_bit_it_2_vnu_181_in_0, msg_to_bit_it_2_vnu_181_in_1, msg_to_bit_it_2_vnu_181_in_2, data_out[181]);
vnu_h hard_dec182(data_182, msg_to_bit_it_2_vnu_182_in_0, msg_to_bit_it_2_vnu_182_in_1, msg_to_bit_it_2_vnu_182_in_2, data_out[182]);
vnu_h hard_dec183(data_183, msg_to_bit_it_2_vnu_183_in_0, msg_to_bit_it_2_vnu_183_in_1, msg_to_bit_it_2_vnu_183_in_2, data_out[183]);
vnu_h hard_dec184(data_184, msg_to_bit_it_2_vnu_184_in_0, msg_to_bit_it_2_vnu_184_in_1, msg_to_bit_it_2_vnu_184_in_2, data_out[184]);
vnu_h hard_dec185(data_185, msg_to_bit_it_2_vnu_185_in_0, msg_to_bit_it_2_vnu_185_in_1, msg_to_bit_it_2_vnu_185_in_2, data_out[185]);
vnu_h hard_dec186(data_186, msg_to_bit_it_2_vnu_186_in_0, msg_to_bit_it_2_vnu_186_in_1, msg_to_bit_it_2_vnu_186_in_2, data_out[186]);
vnu_h hard_dec187(data_187, msg_to_bit_it_2_vnu_187_in_0, msg_to_bit_it_2_vnu_187_in_1, msg_to_bit_it_2_vnu_187_in_2, data_out[187]);
vnu_h hard_dec188(data_188, msg_to_bit_it_2_vnu_188_in_0, msg_to_bit_it_2_vnu_188_in_1, msg_to_bit_it_2_vnu_188_in_2, data_out[188]);
vnu_h hard_dec189(data_189, msg_to_bit_it_2_vnu_189_in_0, msg_to_bit_it_2_vnu_189_in_1, msg_to_bit_it_2_vnu_189_in_2, data_out[189]);
vnu_h hard_dec190(data_190, msg_to_bit_it_2_vnu_190_in_0, msg_to_bit_it_2_vnu_190_in_1, msg_to_bit_it_2_vnu_190_in_2, data_out[190]);
vnu_h hard_dec191(data_191, msg_to_bit_it_2_vnu_191_in_0, msg_to_bit_it_2_vnu_191_in_1, msg_to_bit_it_2_vnu_191_in_2, data_out[191]);
vnu_h hard_dec192(data_192, msg_to_bit_it_2_vnu_192_in_0, msg_to_bit_it_2_vnu_192_in_1, msg_to_bit_it_2_vnu_192_in_2, data_out[192]);
vnu_h hard_dec193(data_193, msg_to_bit_it_2_vnu_193_in_0, msg_to_bit_it_2_vnu_193_in_1, msg_to_bit_it_2_vnu_193_in_2, data_out[193]);
vnu_h hard_dec194(data_194, msg_to_bit_it_2_vnu_194_in_0, msg_to_bit_it_2_vnu_194_in_1, msg_to_bit_it_2_vnu_194_in_2, data_out[194]);
vnu_h hard_dec195(data_195, msg_to_bit_it_2_vnu_195_in_0, msg_to_bit_it_2_vnu_195_in_1, msg_to_bit_it_2_vnu_195_in_2, data_out[195]);
vnu_h hard_dec196(data_196, msg_to_bit_it_2_vnu_196_in_0, msg_to_bit_it_2_vnu_196_in_1, msg_to_bit_it_2_vnu_196_in_2, data_out[196]);
vnu_h hard_dec197(data_197, msg_to_bit_it_2_vnu_197_in_0, msg_to_bit_it_2_vnu_197_in_1, msg_to_bit_it_2_vnu_197_in_2, data_out[197]);



//perform hard decision decoding


endmodule